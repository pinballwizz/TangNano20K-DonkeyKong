library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity dkong_wav is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of dkong_wav is
	type rom is array(0 to  39167) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7D",X"7D",X"7D",X"7D",X"7C",X"7A",X"6D",X"4D",X"37",X"34",X"40",
		X"52",X"7F",X"AD",X"BD",X"C2",X"BF",X"B7",X"B0",X"A7",X"9E",X"8F",X"6A",X"4D",X"41",X"46",X"52",
		X"77",X"A5",X"B9",X"BD",X"B9",X"B1",X"A8",X"A1",X"98",X"8F",X"76",X"53",X"3E",X"3B",X"41",X"58",
		X"87",X"A7",X"B1",X"B1",X"AD",X"A5",X"9E",X"96",X"8D",X"86",X"6B",X"4C",X"3B",X"3A",X"43",X"5B",
		X"87",X"A4",X"AD",X"AD",X"A7",X"A1",X"99",X"93",X"8C",X"84",X"6E",X"50",X"3E",X"3B",X"41",X"55",
		X"80",X"9F",X"A8",X"AB",X"A5",X"9F",X"99",X"93",X"8D",X"87",X"7C",X"5F",X"47",X"3E",X"41",X"4C",
		X"6A",X"92",X"A4",X"AA",X"A7",X"A2",X"9C",X"95",X"90",X"8A",X"84",X"76",X"59",X"46",X"41",X"47",
		X"55",X"77",X"98",X"A4",X"A8",X"A5",X"9F",X"99",X"93",X"8F",X"89",X"84",X"76",X"5B",X"49",X"46",
		X"4A",X"58",X"79",X"98",X"A4",X"A7",X"A4",X"9F",X"99",X"93",X"8F",X"89",X"84",X"79",X"61",X"4F",
		X"49",X"4C",X"56",X"71",X"92",X"A1",X"A4",X"A2",X"9E",X"98",X"93",X"8F",X"8A",X"86",X"7F",X"6A",
		X"56",X"4C",X"4D",X"55",X"68",X"89",X"9B",X"A2",X"A2",X"9F",X"99",X"95",X"90",X"8C",X"87",X"83",
		X"76",X"61",X"52",X"4F",X"53",X"5E",X"7A",X"93",X"9E",X"A2",X"9F",X"9B",X"96",X"92",X"8D",X"89",
		X"84",X"80",X"6E",X"5B",X"52",X"52",X"58",X"67",X"84",X"98",X"9F",X"9F",X"9C",X"98",X"93",X"90",
		X"8C",X"87",X"83",X"7D",X"6B",X"5B",X"53",X"55",X"5B",X"6D",X"87",X"98",X"9C",X"9C",X"99",X"95",
		X"90",X"8D",X"89",X"86",X"83",X"7C",X"6B",X"5C",X"56",X"58",X"5E",X"6E",X"89",X"96",X"9B",X"9B",
		X"99",X"95",X"90",X"8C",X"89",X"86",X"83",X"7D",X"6E",X"5F",X"59",X"59",X"5F",X"6D",X"84",X"93",
		X"99",X"9B",X"98",X"93",X"90",X"8C",X"89",X"86",X"83",X"7F",X"71",X"64",X"5C",X"5B",X"5F",X"6B",
		X"81",X"90",X"98",X"98",X"96",X"93",X"8F",X"8C",X"89",X"86",X"83",X"80",X"77",X"68",X"5F",X"5E",
		X"61",X"68",X"7C",X"8D",X"95",X"98",X"96",X"93",X"90",X"8C",X"89",X"86",X"84",X"81",X"7C",X"6D",
		X"62",X"5F",X"61",X"65",X"74",X"87",X"92",X"96",X"95",X"92",X"8F",X"8C",X"89",X"87",X"84",X"81",
		X"7F",X"76",X"68",X"62",X"62",X"65",X"6D",X"80",X"8D",X"93",X"95",X"92",X"90",X"8D",X"8A",X"87",
		X"86",X"83",X"80",X"7C",X"70",X"65",X"62",X"64",X"68",X"76",X"87",X"90",X"93",X"92",X"90",X"8D",
		X"8A",X"89",X"86",X"83",X"81",X"7F",X"77",X"6B",X"64",X"64",X"67",X"6D",X"7D",X"8C",X"90",X"93",
		X"92",X"8F",X"8C",X"8A",X"87",X"84",X"83",X"81",X"7D",X"73",X"6A",X"65",X"67",X"6A",X"73",X"83",
		X"8D",X"90",X"90",X"8F",X"8D",X"8A",X"87",X"86",X"84",X"81",X"80",X"7A",X"70",X"68",X"67",X"68",
		X"6D",X"77",X"86",X"8D",X"90",X"8F",X"8D",X"8C",X"89",X"87",X"84",X"83",X"80",X"7F",X"79",X"6E",
		X"6A",X"68",X"6B",X"70",X"7D",X"89",X"8D",X"8F",X"8F",X"8C",X"8A",X"87",X"86",X"84",X"83",X"81",
		X"7F",X"77",X"6E",X"6A",X"6A",X"6D",X"73",X"80",X"8A",X"8D",X"8F",X"8D",X"8C",X"89",X"87",X"84",
		X"83",X"81",X"80",X"7D",X"76",X"6E",X"6B",X"6B",X"6E",X"76",X"81",X"8A",X"8D",X"8D",X"8C",X"8A",
		X"87",X"86",X"84",X"83",X"81",X"80",X"7D",X"74",X"6E",X"6D",X"6D",X"70",X"77",X"83",X"8A",X"8D",
		X"8D",X"8C",X"8A",X"87",X"86",X"84",X"83",X"81",X"80",X"7C",X"74",X"6E",X"6D",X"6E",X"71",X"79",
		X"84",X"8A",X"8C",X"8C",X"8A",X"89",X"87",X"84",X"83",X"81",X"81",X"80",X"7D",X"76",X"70",X"6E",
		X"6E",X"71",X"77",X"81",X"89",X"8C",X"8C",X"8A",X"89",X"87",X"86",X"84",X"83",X"81",X"80",X"80",
		X"7F",X"7C",X"76",X"70",X"6E",X"6E",X"71",X"77",X"81",X"89",X"8A",X"8A",X"8A",X"87",X"86",X"86",
		X"84",X"83",X"81",X"81",X"81",X"80",X"80",X"86",X"92",X"96",X"96",X"93",X"8D",X"81",X"73",X"6A",
		X"65",X"65",X"67",X"6A",X"6D",X"6E",X"71",X"74",X"77",X"79",X"7C",X"7F",X"89",X"93",X"98",X"98",
		X"95",X"8F",X"80",X"73",X"6B",X"68",X"6A",X"6D",X"70",X"73",X"76",X"79",X"7A",X"7D",X"7F",X"81",
		X"8A",X"96",X"9B",X"9B",X"98",X"92",X"84",X"76",X"6E",X"6B",X"6D",X"6E",X"71",X"74",X"77",X"79",
		X"7C",X"7D",X"80",X"83",X"8F",X"99",X"9C",X"9B",X"96",X"8F",X"7F",X"73",X"6D",X"6B",X"6D",X"6E",
		X"73",X"74",X"77",X"7A",X"7C",X"7F",X"81",X"89",X"95",X"9B",X"9B",X"98",X"93",X"84",X"76",X"6E",
		X"6B",X"6D",X"6E",X"71",X"74",X"77",X"7A",X"7C",X"7F",X"80",X"87",X"95",X"9B",X"9B",X"98",X"93",
		X"87",X"77",X"6E",X"6B",X"6D",X"6E",X"71",X"74",X"76",X"79",X"7C",X"7D",X"80",X"87",X"93",X"9B",
		X"9B",X"96",X"92",X"84",X"76",X"6E",X"6B",X"6D",X"6E",X"71",X"74",X"77",X"79",X"7C",X"7D",X"80",
		X"8A",X"96",X"9B",X"99",X"96",X"8F",X"80",X"73",X"6D",X"6B",X"6D",X"70",X"73",X"74",X"77",X"7A",
		X"7C",X"7F",X"83",X"8F",X"98",X"9B",X"98",X"93",X"8A",X"7A",X"70",X"6B",X"6B",X"6D",X"70",X"73",
		X"76",X"77",X"7A",X"7D",X"7F",X"89",X"95",X"99",X"99",X"96",X"8F",X"81",X"73",X"6D",X"6B",X"6D",
		X"70",X"73",X"74",X"77",X"79",X"7C",X"7F",X"84",X"90",X"98",X"99",X"96",X"92",X"86",X"77",X"6E",
		X"6B",X"6D",X"6E",X"71",X"74",X"77",X"79",X"7C",X"7F",X"81",X"8D",X"96",X"99",X"98",X"93",X"8A",
		X"7C",X"71",X"6D",X"6D",X"6E",X"71",X"74",X"76",X"79",X"7A",X"7D",X"80",X"8A",X"95",X"98",X"96",
		X"93",X"8D",X"7F",X"73",X"6E",X"6D",X"6E",X"71",X"74",X"76",X"79",X"7A",X"7D",X"7F",X"87",X"92",
		X"96",X"98",X"95",X"8F",X"81",X"74",X"6E",X"6D",X"6E",X"71",X"74",X"76",X"79",X"7A",X"7D",X"7F",
		X"86",X"90",X"96",X"96",X"93",X"8F",X"83",X"76",X"70",X"6E",X"6E",X"71",X"74",X"76",X"79",X"7A",
		X"7D",X"7F",X"84",X"8F",X"95",X"95",X"93",X"8F",X"83",X"77",X"71",X"70",X"70",X"71",X"74",X"76",
		X"79",X"7A",X"7D",X"7F",X"83",X"8D",X"92",X"93",X"92",X"8F",X"84",X"79",X"73",X"70",X"71",X"73",
		X"76",X"77",X"79",X"7A",X"7C",X"7F",X"83",X"8C",X"92",X"93",X"92",X"8F",X"84",X"7A",X"74",X"71",
		X"71",X"73",X"76",X"77",X"79",X"7A",X"7D",X"7F",X"81",X"8A",X"90",X"92",X"90",X"8D",X"86",X"7A",
		X"74",X"71",X"73",X"74",X"76",X"77",X"7A",X"7A",X"7C",X"7F",X"81",X"89",X"8F",X"90",X"8F",X"8C",
		X"86",X"7C",X"76",X"73",X"73",X"74",X"76",X"79",X"79",X"7A",X"7D",X"7F",X"80",X"87",X"8D",X"8F",
		X"8D",X"8C",X"86",X"7C",X"77",X"74",X"74",X"76",X"77",X"79",X"7A",X"7C",X"7D",X"7D",X"80",X"86",
		X"8C",X"8D",X"8D",X"8C",X"86",X"7F",X"77",X"76",X"74",X"76",X"77",X"79",X"7A",X"7C",X"7C",X"7D",
		X"80",X"84",X"8A",X"8D",X"8C",X"8A",X"86",X"7F",X"79",X"76",X"76",X"76",X"77",X"79",X"7A",X"7C",
		X"7D",X"7F",X"7F",X"83",X"8A",X"8C",X"8C",X"8A",X"87",X"7F",X"79",X"76",X"76",X"77",X"77",X"79",
		X"7A",X"7C",X"7D",X"7F",X"7F",X"84",X"89",X"8A",X"8C",X"8A",X"87",X"80",X"7A",X"77",X"77",X"77",
		X"79",X"7A",X"7A",X"7C",X"7D",X"7F",X"7F",X"83",X"87",X"8A",X"8A",X"89",X"87",X"80",X"7A",X"79",
		X"77",X"79",X"79",X"7A",X"7C",X"7C",X"7D",X"7F",X"7F",X"81",X"86",X"89",X"89",X"89",X"86",X"80",
		X"7C",X"79",X"77",X"79",X"79",X"7A",X"7C",X"7C",X"7D",X"7D",X"7F",X"81",X"86",X"89",X"89",X"89",
		X"87",X"81",X"7C",X"79",X"79",X"79",X"7A",X"7A",X"7C",X"7D",X"7D",X"7F",X"7F",X"81",X"86",X"87",
		X"89",X"87",X"86",X"81",X"7C",X"79",X"79",X"79",X"79",X"7A",X"7C",X"7C",X"7D",X"7F",X"7F",X"81",
		X"86",X"87",X"87",X"87",X"84",X"80",X"7C",X"7A",X"79",X"7A",X"7A",X"7C",X"7C",X"7D",X"7D",X"7F",
		X"83",X"86",X"87",X"86",X"86",X"83",X"7D",X"7A",X"79",X"7A",X"7A",X"7C",X"7C",X"7D",X"7D",X"7F",
		X"83",X"86",X"86",X"86",X"84",X"81",X"7D",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7D",X"7F",X"81",
		X"84",X"86",X"86",X"84",X"83",X"7F",X"7C",X"7A",X"7A",X"7A",X"7C",X"7D",X"7D",X"7F",X"81",X"84",
		X"86",X"84",X"83",X"81",X"7D",X"7A",X"7A",X"7A",X"7A",X"7C",X"7D",X"7D",X"80",X"83",X"84",X"84",
		X"84",X"83",X"7F",X"7C",X"7A",X"7A",X"7C",X"7C",X"7D",X"7D",X"80",X"83",X"84",X"84",X"84",X"83",
		X"7F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7F",X"80",X"83",X"84",X"84",X"84",X"81",X"7F",X"7C",
		X"7C",X"7C",X"7C",X"7D",X"7D",X"7F",X"81",X"83",X"84",X"84",X"83",X"80",X"7D",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7F",X"80",X"83",X"84",X"84",X"83",X"81",X"7F",X"7D",X"7C",X"7C",X"7D",X"7D",X"7F",
		X"80",X"81",X"83",X"83",X"83",X"81",X"7F",X"7D",X"7C",X"7C",X"7C",X"7D",X"7D",X"80",X"81",X"83",
		X"83",X"83",X"81",X"7F",X"7D",X"7C",X"7C",X"7C",X"7D",X"7D",X"80",X"81",X"81",X"83",X"83",X"81",
		X"7F",X"7D",X"7C",X"7C",X"7C",X"7D",X"7F",X"80",X"83",X"83",X"83",X"83",X"81",X"7F",X"7D",X"7C",
		X"7C",X"7D",X"7D",X"7F",X"80",X"81",X"83",X"83",X"81",X"80",X"7D",X"7C",X"7C",X"7C",X"7D",X"7D",
		X"80",X"81",X"81",X"83",X"81",X"81",X"7F",X"7D",X"7C",X"7D",X"7D",X"7D",X"7F",X"80",X"81",X"83",
		X"83",X"81",X"80",X"7F",X"7D",X"7D",X"7C",X"7D",X"7D",X"7F",X"80",X"81",X"83",X"81",X"81",X"7F",
		X"7D",X"7D",X"7C",X"7D",X"7D",X"7F",X"80",X"81",X"81",X"81",X"81",X"80",X"7F",X"7D",X"7D",X"7D",
		X"7D",X"7F",X"80",X"81",X"81",X"81",X"81",X"81",X"7F",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"80",
		X"81",X"81",X"81",X"81",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"80",X"81",X"81",X"81",X"81",
		X"80",X"7F",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"80",X"81",X"81",X"81",X"80",X"7F",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7F",X"80",X"81",X"81",X"81",X"81",X"80",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",
		X"80",X"81",X"81",X"81",X"81",X"80",X"7F",X"7D",X"7D",X"7F",X"7F",X"7F",X"80",X"81",X"81",X"81",
		X"81",X"80",X"7F",X"7D",X"7D",X"7D",X"7D",X"7F",X"80",X"80",X"81",X"81",X"81",X"80",X"7F",X"7D",
		X"7D",X"7D",X"7D",X"7F",X"80",X"81",X"81",X"81",X"81",X"80",X"7F",X"7D",X"7D",X"7D",X"7D",X"7F",
		X"7F",X"80",X"81",X"81",X"81",X"80",X"7F",X"7F",X"7D",X"7D",X"7F",X"7F",X"7F",X"80",X"80",X"81",
		X"81",X"80",X"80",X"7F",X"7D",X"7D",X"7D",X"7F",X"7F",X"80",X"80",X"81",X"81",X"80",X"80",X"7F",
		X"7D",X"7D",X"7D",X"7F",X"7F",X"80",X"80",X"81",X"81",X"80",X"80",X"7F",X"7D",X"7D",X"7D",X"7D",
		X"7F",X"80",X"80",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7D",X"7D",X"7F",X"7F",X"80",X"80",X"80",
		X"81",X"81",X"80",X"7F",X"7F",X"7D",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",X"80",X"80",X"7F",
		X"7F",X"7D",X"7D",X"7F",X"7F",X"80",X"80",X"80",X"80",X"81",X"80",X"7F",X"7D",X"7D",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"81",X"80",X"80",X"80",X"7F",X"7D",X"7D",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"80",X"80",X"80",
		X"7F",X"7D",X"7F",X"7D",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"7D",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",
		X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",
		X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"7C",X"7C",X"7C",X"7A",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7E",X"7E",X"7E",X"80",X"7E",X"7E",X"7E",X"7E",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7C",X"7E",X"80",X"82",X"84",X"86",X"84",X"84",X"82",X"82",X"7C",X"7A",X"78",
		X"76",X"76",X"76",X"76",X"78",X"78",X"7A",X"7C",X"7C",X"7E",X"84",X"88",X"8C",X"8E",X"8C",X"8C",
		X"8A",X"88",X"80",X"7A",X"74",X"72",X"72",X"72",X"72",X"74",X"76",X"78",X"78",X"7A",X"7C",X"80",
		X"88",X"8E",X"94",X"96",X"96",X"94",X"92",X"8E",X"84",X"7A",X"72",X"6E",X"6C",X"6C",X"6E",X"6E",
		X"70",X"72",X"76",X"78",X"7A",X"7C",X"82",X"8A",X"92",X"98",X"9A",X"9C",X"9C",X"9A",X"94",X"88",
		X"7A",X"70",X"6C",X"68",X"68",X"6A",X"6A",X"6E",X"70",X"74",X"76",X"7A",X"7C",X"7E",X"84",X"8E",
		X"94",X"9A",X"9C",X"9E",X"9E",X"9C",X"96",X"84",X"76",X"6E",X"68",X"64",X"66",X"66",X"6A",X"6C",
		X"70",X"72",X"76",X"78",X"7C",X"7E",X"82",X"88",X"90",X"96",X"9C",X"9E",X"A0",X"A0",X"9E",X"94",
		X"84",X"76",X"6C",X"66",X"64",X"64",X"66",X"68",X"6A",X"6E",X"70",X"74",X"76",X"7A",X"7E",X"80",
		X"84",X"8A",X"92",X"98",X"9E",X"A0",X"A0",X"A0",X"9C",X"8E",X"7C",X"70",X"68",X"64",X"64",X"64",
		X"66",X"68",X"6C",X"6E",X"72",X"74",X"78",X"7A",X"7E",X"80",X"82",X"86",X"8E",X"96",X"9C",X"9E",
		X"A0",X"A0",X"A0",X"9A",X"8A",X"78",X"6E",X"68",X"64",X"62",X"64",X"66",X"6A",X"6C",X"6E",X"72",
		X"74",X"78",X"7A",X"7E",X"80",X"82",X"84",X"8C",X"94",X"9A",X"9C",X"A0",X"A0",X"A0",X"9E",X"94",
		X"80",X"74",X"6A",X"64",X"62",X"64",X"66",X"68",X"6A",X"6E",X"70",X"72",X"76",X"78",X"7A",X"7C",
		X"7E",X"80",X"82",X"86",X"8E",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9C",X"8C",X"7C",X"70",X"68",
		X"64",X"62",X"64",X"66",X"68",X"6A",X"6E",X"70",X"74",X"76",X"7A",X"7C",X"7E",X"80",X"82",X"82",
		X"84",X"88",X"90",X"98",X"9C",X"A0",X"A0",X"A2",X"A0",X"98",X"88",X"78",X"6C",X"66",X"62",X"62",
		X"64",X"66",X"68",X"6C",X"6E",X"70",X"74",X"76",X"78",X"7C",X"7C",X"7E",X"80",X"82",X"84",X"86",
		X"8E",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9E",X"92",X"80",X"72",X"68",X"64",X"62",X"62",X"64",
		X"66",X"68",X"6C",X"70",X"72",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"82",X"84",X"86",X"88",
		X"90",X"96",X"9C",X"9E",X"A0",X"A0",X"A0",X"9A",X"8A",X"7A",X"6C",X"64",X"62",X"60",X"62",X"64",
		X"66",X"6A",X"6C",X"70",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"82",X"84",X"86",X"86",
		X"8C",X"92",X"98",X"9C",X"A0",X"A2",X"A0",X"A0",X"98",X"86",X"74",X"6A",X"64",X"60",X"60",X"62",
		X"64",X"66",X"6A",X"6C",X"70",X"74",X"76",X"7A",X"7C",X"7E",X"7E",X"80",X"82",X"84",X"84",X"86",
		X"86",X"88",X"8E",X"96",X"9A",X"9E",X"A0",X"A2",X"A0",X"9C",X"92",X"7E",X"70",X"68",X"62",X"60",
		X"60",X"62",X"64",X"68",X"6C",X"70",X"72",X"74",X"78",X"7A",X"7C",X"7E",X"80",X"80",X"82",X"82",
		X"84",X"84",X"86",X"86",X"8A",X"92",X"98",X"9C",X"9E",X"A0",X"A0",X"9E",X"9A",X"8C",X"7A",X"6E",
		X"66",X"62",X"60",X"62",X"64",X"66",X"68",X"6C",X"70",X"72",X"74",X"78",X"7A",X"7C",X"7E",X"80",
		X"82",X"82",X"82",X"84",X"84",X"84",X"86",X"86",X"8C",X"94",X"9A",X"9E",X"9E",X"A0",X"A0",X"9E",
		X"98",X"86",X"74",X"68",X"62",X"60",X"60",X"62",X"64",X"66",X"6A",X"6E",X"70",X"74",X"76",X"78",
		X"7A",X"7C",X"7E",X"80",X"80",X"80",X"82",X"84",X"84",X"86",X"86",X"8C",X"94",X"98",X"9C",X"9E",
		X"A0",X"A0",X"9E",X"9A",X"8A",X"78",X"6C",X"64",X"60",X"60",X"60",X"62",X"66",X"68",X"6C",X"6E",
		X"72",X"74",X"78",X"7A",X"7C",X"7E",X"7E",X"80",X"82",X"82",X"84",X"84",X"84",X"88",X"90",X"98",
		X"9C",X"9E",X"A0",X"A2",X"A0",X"9E",X"92",X"7E",X"70",X"66",X"62",X"60",X"60",X"62",X"64",X"68",
		X"6C",X"6E",X"70",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"82",X"84",X"84",X"86",X"8C",
		X"94",X"9A",X"9E",X"A0",X"A0",X"A0",X"A0",X"9A",X"88",X"78",X"6C",X"64",X"60",X"60",X"62",X"64",
		X"66",X"6A",X"6E",X"70",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"82",X"84",X"86",X"88",
		X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"A0",X"98",X"86",X"76",X"6A",X"64",X"60",X"60",X"62",
		X"64",X"66",X"6A",X"6C",X"70",X"72",X"76",X"7A",X"7C",X"7E",X"7E",X"80",X"82",X"82",X"84",X"86",
		X"88",X"90",X"96",X"9C",X"9E",X"A2",X"A2",X"A0",X"9E",X"92",X"80",X"70",X"68",X"62",X"60",X"62",
		X"62",X"64",X"68",X"6C",X"6E",X"72",X"74",X"76",X"7A",X"7C",X"7E",X"80",X"82",X"84",X"84",X"86",
		X"8A",X"90",X"96",X"9C",X"A0",X"A0",X"A2",X"A0",X"9E",X"90",X"7E",X"70",X"68",X"64",X"62",X"62",
		X"64",X"66",X"6A",X"6C",X"70",X"72",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"80",X"82",X"84",X"86",
		X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9E",X"96",X"84",X"74",X"6A",X"64",X"60",X"60",X"62",
		X"64",X"68",X"6A",X"6E",X"70",X"74",X"76",X"7A",X"7C",X"7E",X"80",X"82",X"82",X"84",X"88",X"90",
		X"96",X"9C",X"A0",X"A2",X"A2",X"A0",X"9E",X"92",X"7E",X"70",X"66",X"62",X"60",X"60",X"62",X"66",
		X"68",X"6C",X"70",X"72",X"76",X"78",X"7A",X"7E",X"7E",X"82",X"82",X"88",X"90",X"98",X"9C",X"A0",
		X"A2",X"A2",X"A0",X"9C",X"8C",X"7A",X"6E",X"66",X"62",X"60",X"62",X"64",X"68",X"6A",X"6E",X"70",
		X"74",X"76",X"7A",X"7C",X"7E",X"82",X"84",X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9E",X"94",
		X"80",X"72",X"68",X"64",X"62",X"62",X"64",X"66",X"6A",X"6C",X"70",X"72",X"76",X"7A",X"7C",X"7E",
		X"82",X"88",X"90",X"98",X"9C",X"A0",X"A2",X"A2",X"A0",X"9C",X"8A",X"78",X"6C",X"66",X"64",X"62",
		X"64",X"66",X"68",X"6C",X"6E",X"72",X"74",X"78",X"7A",X"7E",X"82",X"8A",X"94",X"98",X"9E",X"A0",
		X"A2",X"A2",X"9E",X"94",X"80",X"72",X"6A",X"64",X"62",X"64",X"64",X"68",X"6A",X"6E",X"72",X"74",
		X"78",X"7C",X"7E",X"84",X"8C",X"94",X"9A",X"9E",X"A0",X"A0",X"A0",X"9C",X"8E",X"7C",X"6E",X"66",
		X"64",X"62",X"62",X"64",X"68",X"6C",X"6E",X"72",X"76",X"78",X"7C",X"80",X"8A",X"92",X"98",X"9C",
		X"A0",X"A0",X"A0",X"9C",X"90",X"7C",X"6E",X"68",X"62",X"62",X"64",X"66",X"68",X"6C",X"6E",X"72",
		X"76",X"7A",X"7E",X"84",X"8E",X"94",X"9A",X"9E",X"A0",X"A0",X"A0",X"98",X"86",X"76",X"6C",X"64",
		X"62",X"62",X"64",X"66",X"6A",X"6E",X"70",X"74",X"78",X"7C",X"82",X"8C",X"94",X"9A",X"9E",X"A0",
		X"A0",X"A0",X"98",X"86",X"76",X"6C",X"66",X"64",X"62",X"64",X"68",X"6A",X"6E",X"72",X"76",X"78",
		X"7E",X"86",X"90",X"96",X"9C",X"9E",X"A0",X"A0",X"9E",X"90",X"7E",X"70",X"68",X"64",X"64",X"64",
		X"66",X"68",X"6C",X"70",X"74",X"78",X"7C",X"84",X"8E",X"96",X"9C",X"9E",X"A0",X"A0",X"9E",X"92",
		X"80",X"72",X"68",X"64",X"64",X"64",X"66",X"6A",X"6C",X"70",X"74",X"78",X"7C",X"86",X"90",X"96",
		X"9C",X"9E",X"A0",X"A0",X"9E",X"8E",X"7C",X"6E",X"66",X"64",X"62",X"64",X"66",X"68",X"6C",X"70",
		X"74",X"7A",X"82",X"8E",X"96",X"9A",X"9E",X"A0",X"A0",X"9E",X"94",X"82",X"74",X"6A",X"66",X"64",
		X"64",X"66",X"68",X"6C",X"70",X"74",X"78",X"80",X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"9E",X"96",
		X"84",X"74",X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"78",X"80",X"8A",X"92",X"98",
		X"9C",X"A0",X"A0",X"9E",X"94",X"80",X"72",X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",
		X"7A",X"84",X"8E",X"94",X"9A",X"9E",X"9E",X"9E",X"9C",X"8C",X"7C",X"6E",X"66",X"64",X"64",X"64",
		X"68",X"6C",X"6E",X"72",X"76",X"80",X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"9E",X"92",X"80",X"72",
		X"6A",X"66",X"64",X"66",X"68",X"6A",X"6E",X"72",X"76",X"7E",X"88",X"90",X"98",X"9A",X"9E",X"9E",
		X"9E",X"96",X"84",X"74",X"6C",X"66",X"64",X"64",X"66",X"6A",X"6C",X"70",X"74",X"7C",X"86",X"90",
		X"96",X"9C",X"9E",X"9E",X"9E",X"96",X"84",X"74",X"6A",X"66",X"64",X"64",X"66",X"6A",X"6C",X"70",
		X"76",X"7E",X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"9E",X"94",X"80",X"72",X"6A",X"66",X"64",X"66",
		X"68",X"6A",X"6E",X"72",X"78",X"82",X"8C",X"92",X"9A",X"9E",X"9E",X"9E",X"9C",X"8C",X"7A",X"6E",
		X"66",X"62",X"62",X"64",X"68",X"6C",X"70",X"74",X"7C",X"88",X"90",X"98",X"9C",X"9E",X"9E",X"9E",
		X"96",X"84",X"74",X"6A",X"66",X"64",X"66",X"66",X"6A",X"6E",X"72",X"78",X"82",X"8C",X"94",X"98",
		X"9C",X"9E",X"9E",X"9A",X"8A",X"78",X"6E",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"80",
		X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"9C",X"8E",X"7C",X"70",X"68",X"64",X"64",X"66",X"68",X"6C",
		X"6E",X"74",X"7C",X"88",X"90",X"96",X"9A",X"9E",X"9E",X"9C",X"90",X"7E",X"72",X"68",X"66",X"64",
		X"66",X"68",X"6C",X"6E",X"72",X"7C",X"86",X"90",X"96",X"9A",X"9C",X"9E",X"9C",X"92",X"7E",X"72",
		X"68",X"64",X"64",X"64",X"68",X"6A",X"6E",X"74",X"7E",X"88",X"90",X"96",X"9A",X"9E",X"9E",X"9C",
		X"90",X"7C",X"70",X"6A",X"66",X"64",X"66",X"68",X"6C",X"6E",X"74",X"7E",X"8A",X"92",X"96",X"9C",
		X"9E",X"9E",X"9C",X"8E",X"7C",X"70",X"68",X"64",X"64",X"66",X"68",X"6C",X"70",X"76",X"80",X"8A",
		X"92",X"98",X"9C",X"9E",X"9E",X"9A",X"88",X"78",X"6E",X"66",X"64",X"64",X"66",X"6A",X"6E",X"72",
		X"7A",X"86",X"8E",X"94",X"9A",X"9C",X"9E",X"9E",X"96",X"84",X"74",X"6A",X"66",X"64",X"64",X"66",
		X"68",X"6C",X"72",X"7C",X"88",X"90",X"96",X"9A",X"9E",X"9E",X"9C",X"90",X"7E",X"70",X"68",X"66",
		X"64",X"66",X"68",X"6C",X"70",X"78",X"82",X"8C",X"94",X"98",X"9C",X"9E",X"9E",X"9A",X"88",X"78",
		X"6C",X"66",X"64",X"64",X"66",X"6A",X"6E",X"72",X"7C",X"86",X"90",X"96",X"9A",X"9E",X"9E",X"9C",
		X"90",X"7E",X"70",X"68",X"64",X"64",X"64",X"68",X"6C",X"6E",X"76",X"82",X"8A",X"94",X"98",X"9C",
		X"9E",X"9E",X"98",X"86",X"74",X"6A",X"66",X"62",X"64",X"66",X"6A",X"6C",X"72",X"7E",X"88",X"90",
		X"96",X"9C",X"9E",X"9E",X"9A",X"8C",X"7A",X"70",X"68",X"64",X"64",X"66",X"68",X"6C",X"72",X"7A",
		X"86",X"8E",X"94",X"9A",X"9E",X"9E",X"9C",X"92",X"7E",X"72",X"68",X"64",X"64",X"66",X"68",X"6C",
		X"6E",X"76",X"82",X"8C",X"94",X"98",X"9C",X"9E",X"9E",X"96",X"82",X"74",X"6C",X"66",X"64",X"66",
		X"68",X"6A",X"6E",X"72",X"7C",X"86",X"90",X"96",X"9A",X"9E",X"9E",X"9E",X"92",X"80",X"72",X"6A",
		X"66",X"64",X"66",X"68",X"6A",X"6E",X"72",X"7A",X"86",X"8E",X"96",X"9A",X"9E",X"A0",X"9E",X"94",
		X"82",X"74",X"6C",X"66",X"64",X"66",X"68",X"6A",X"6E",X"72",X"78",X"80",X"8A",X"94",X"98",X"9C",
		X"9E",X"A0",X"9C",X"8C",X"7A",X"6E",X"68",X"64",X"64",X"64",X"68",X"6C",X"6E",X"72",X"7A",X"82",
		X"8C",X"94",X"9A",X"9E",X"A0",X"A0",X"9C",X"8C",X"7A",X"6E",X"68",X"64",X"64",X"66",X"68",X"6C",
		X"70",X"74",X"78",X"80",X"8A",X"92",X"9A",X"9C",X"9E",X"9E",X"9C",X"92",X"7E",X"72",X"68",X"64",
		X"64",X"66",X"68",X"6A",X"6E",X"70",X"74",X"7A",X"84",X"8E",X"94",X"9A",X"9E",X"9E",X"9E",X"9C",
		X"8C",X"7A",X"6E",X"68",X"64",X"64",X"66",X"68",X"6A",X"6E",X"72",X"76",X"7A",X"84",X"8E",X"96",
		X"9A",X"9E",X"A0",X"9E",X"9C",X"8C",X"7C",X"6E",X"68",X"66",X"64",X"66",X"68",X"6A",X"6E",X"72",
		X"76",X"78",X"80",X"8A",X"92",X"9A",X"9C",X"A0",X"A0",X"A0",X"96",X"82",X"74",X"6A",X"66",X"64",
		X"64",X"66",X"68",X"6C",X"70",X"72",X"76",X"7C",X"84",X"8E",X"94",X"9A",X"9E",X"A0",X"A0",X"9E",
		X"92",X"80",X"72",X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"76",X"7A",X"82",X"8E",
		X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"94",X"82",X"74",X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",
		X"70",X"72",X"76",X"7A",X"7E",X"88",X"92",X"98",X"9E",X"A0",X"A0",X"A0",X"9C",X"8C",X"7A",X"6E",
		X"68",X"64",X"64",X"66",X"66",X"6A",X"6C",X"70",X"72",X"78",X"7A",X"80",X"88",X"92",X"9A",X"9C",
		X"A0",X"A0",X"A0",X"9C",X"8A",X"7A",X"6E",X"68",X"64",X"64",X"66",X"68",X"6A",X"6E",X"72",X"74",
		X"78",X"7C",X"80",X"88",X"92",X"98",X"9C",X"A0",X"A0",X"A0",X"9E",X"90",X"7C",X"70",X"68",X"64",
		X"64",X"64",X"66",X"68",X"6C",X"6E",X"72",X"76",X"78",X"7E",X"84",X"8E",X"96",X"9A",X"9E",X"A0",
		X"A0",X"9E",X"96",X"84",X"74",X"6C",X"66",X"64",X"64",X"66",X"68",X"6A",X"6E",X"72",X"74",X"78",
		X"7C",X"80",X"88",X"90",X"98",X"9C",X"9E",X"A0",X"A0",X"A0",X"94",X"80",X"72",X"6A",X"64",X"64",
		X"64",X"66",X"68",X"6C",X"6E",X"72",X"74",X"78",X"7C",X"7E",X"88",X"90",X"98",X"9C",X"9E",X"A0",
		X"A0",X"9E",X"94",X"82",X"72",X"6A",X"64",X"62",X"64",X"64",X"68",X"6A",X"6E",X"70",X"74",X"78",
		X"7A",X"7E",X"84",X"8E",X"94",X"9A",X"9E",X"A0",X"A0",X"A0",X"9A",X"8A",X"78",X"6C",X"66",X"64",
		X"62",X"64",X"66",X"6A",X"6C",X"70",X"72",X"76",X"7A",X"7C",X"80",X"88",X"90",X"98",X"9C",X"A0",
		X"A2",X"A0",X"A0",X"96",X"84",X"74",X"6A",X"64",X"62",X"64",X"64",X"68",X"6A",X"6E",X"70",X"74",
		X"78",X"7A",X"7E",X"82",X"8A",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9E",X"92",X"7E",X"70",X"68",
		X"62",X"62",X"64",X"64",X"68",X"6C",X"6E",X"72",X"76",X"7A",X"7C",X"80",X"84",X"8C",X"94",X"9A",
		X"9E",X"A0",X"A2",X"A0",X"9E",X"92",X"7E",X"72",X"6A",X"64",X"62",X"64",X"66",X"68",X"6A",X"6E",
		X"70",X"74",X"78",X"7A",X"7E",X"80",X"88",X"90",X"96",X"9C",X"9E",X"A0",X"A0",X"9E",X"96",X"84",
		X"74",X"6A",X"64",X"62",X"62",X"64",X"66",X"6A",X"6E",X"70",X"74",X"76",X"7A",X"7C",X"7E",X"84",
		X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A2",X"9E",X"8E",X"7C",X"70",X"68",X"64",X"62",X"64",X"64",
		X"68",X"6A",X"6E",X"72",X"74",X"78",X"7A",X"7E",X"80",X"88",X"90",X"96",X"9C",X"A0",X"A2",X"A2",
		X"A2",X"98",X"86",X"76",X"6A",X"66",X"62",X"62",X"64",X"66",X"6A",X"6C",X"70",X"72",X"76",X"78",
		X"7C",X"7E",X"82",X"8A",X"92",X"98",X"9E",X"A0",X"A2",X"A2",X"A0",X"96",X"82",X"74",X"6A",X"64",
		X"62",X"62",X"64",X"68",X"6A",X"6E",X"70",X"74",X"76",X"78",X"7C",X"7E",X"82",X"8A",X"92",X"9A",
		X"9E",X"A0",X"A2",X"A0",X"9E",X"94",X"80",X"72",X"6A",X"64",X"62",X"64",X"64",X"68",X"6A",X"6E",
		X"70",X"74",X"76",X"7A",X"7C",X"7E",X"82",X"8A",X"92",X"98",X"9E",X"A0",X"A2",X"A2",X"A0",X"96",
		X"82",X"74",X"6A",X"64",X"62",X"62",X"62",X"66",X"6A",X"6C",X"70",X"74",X"76",X"7A",X"7C",X"80",
		X"82",X"8A",X"92",X"98",X"9E",X"A0",X"A2",X"A0",X"A0",X"9A",X"88",X"78",X"6C",X"66",X"62",X"62",
		X"64",X"66",X"6A",X"6C",X"70",X"72",X"76",X"78",X"7C",X"7E",X"80",X"84",X"8C",X"94",X"9A",X"9E",
		X"A0",X"A2",X"A0",X"9C",X"8E",X"7C",X"70",X"66",X"62",X"62",X"62",X"64",X"66",X"6A",X"6E",X"70",
		X"74",X"76",X"7A",X"7C",X"80",X"82",X"8A",X"92",X"98",X"9E",X"A0",X"A2",X"A2",X"A0",X"98",X"86",
		X"76",X"6A",X"64",X"62",X"62",X"64",X"66",X"6A",X"6C",X"6E",X"72",X"74",X"78",X"7C",X"7E",X"80",
		X"84",X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9E",X"92",X"80",X"72",X"68",X"64",X"62",X"62",
		X"64",X"66",X"6A",X"6E",X"70",X"74",X"76",X"78",X"7C",X"7E",X"80",X"86",X"8E",X"96",X"9A",X"9E",
		X"A0",X"A2",X"A2",X"9C",X"8C",X"7C",X"6E",X"66",X"64",X"62",X"64",X"64",X"68",X"6A",X"6E",X"70",
		X"74",X"78",X"7A",X"7E",X"80",X"82",X"88",X"92",X"98",X"9C",X"A0",X"A2",X"A0",X"A0",X"9A",X"88",
		X"78",X"6C",X"64",X"62",X"60",X"62",X"64",X"68",X"6A",X"6E",X"72",X"76",X"78",X"7C",X"80",X"82",
		X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9E",X"92",X"80",X"70",X"68",X"62",X"62",X"62",X"64",
		X"66",X"6A",X"6E",X"72",X"74",X"78",X"7C",X"7E",X"84",X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",
		X"9E",X"90",X"7C",X"70",X"68",X"64",X"62",X"62",X"66",X"68",X"6C",X"6E",X"72",X"74",X"78",X"7C",
		X"80",X"8A",X"92",X"98",X"9E",X"A0",X"A2",X"A0",X"9E",X"90",X"7E",X"70",X"68",X"64",X"62",X"62",
		X"64",X"68",X"6A",X"6E",X"72",X"74",X"78",X"7C",X"82",X"8C",X"94",X"9A",X"9E",X"A0",X"A0",X"A0",
		X"9A",X"88",X"78",X"6C",X"66",X"64",X"62",X"66",X"68",X"6A",X"6E",X"70",X"74",X"78",X"7A",X"82",
		X"8C",X"94",X"9A",X"9E",X"A0",X"A0",X"A0",X"9A",X"86",X"76",X"6C",X"66",X"62",X"62",X"64",X"66",
		X"6A",X"6E",X"70",X"74",X"78",X"7E",X"86",X"90",X"96",X"9C",X"9E",X"A0",X"A0",X"9E",X"92",X"7E",
		X"70",X"68",X"64",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"76",X"7C",X"86",X"8E",X"96",X"9C",
		X"9E",X"A0",X"A0",X"9E",X"92",X"80",X"72",X"6A",X"64",X"62",X"64",X"66",X"68",X"6C",X"70",X"74",
		X"76",X"7C",X"86",X"90",X"96",X"9C",X"A0",X"A0",X"A0",X"9E",X"90",X"7C",X"70",X"68",X"64",X"64",
		X"64",X"66",X"6A",X"6C",X"70",X"74",X"78",X"80",X"8C",X"94",X"9A",X"9C",X"A0",X"A0",X"A0",X"96",
		X"84",X"74",X"6C",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"78",X"7E",X"8A",X"92",X"98",
		X"9C",X"A0",X"A0",X"A0",X"98",X"88",X"76",X"6C",X"66",X"64",X"64",X"66",X"68",X"6C",X"6E",X"72",
		X"76",X"80",X"8A",X"92",X"98",X"9C",X"9E",X"A0",X"9E",X"96",X"84",X"76",X"6A",X"64",X"62",X"62",
		X"66",X"68",X"6C",X"70",X"72",X"78",X"82",X"8C",X"94",X"98",X"9C",X"9E",X"9E",X"9E",X"92",X"80",
		X"72",X"68",X"64",X"64",X"64",X"66",X"6A",X"6E",X"70",X"74",X"7C",X"86",X"90",X"96",X"9A",X"9E",
		X"9E",X"A0",X"98",X"86",X"76",X"6C",X"66",X"64",X"64",X"66",X"6A",X"6C",X"70",X"74",X"7A",X"84",
		X"8E",X"94",X"9A",X"9E",X"9E",X"9E",X"9A",X"8A",X"7A",X"6E",X"66",X"64",X"64",X"66",X"68",X"6C",
		X"6E",X"72",X"78",X"82",X"8C",X"94",X"9A",X"9C",X"A0",X"A0",X"9C",X"8A",X"7A",X"6E",X"66",X"64",
		X"64",X"66",X"68",X"6C",X"6E",X"74",X"7A",X"86",X"8E",X"96",X"9A",X"9E",X"A0",X"A0",X"9A",X"88",
		X"78",X"6C",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"7C",X"88",X"90",X"98",X"9C",X"9E",
		X"A0",X"9E",X"94",X"82",X"74",X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"76",X"82",X"8C",
		X"94",X"9A",X"9E",X"A0",X"A0",X"9A",X"8A",X"7A",X"6E",X"68",X"64",X"64",X"66",X"68",X"6C",X"70",
		X"74",X"7E",X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"9C",X"92",X"7E",X"70",X"68",X"64",X"64",X"64",
		X"68",X"6A",X"6E",X"72",X"7A",X"86",X"8E",X"96",X"9A",X"9E",X"A0",X"9E",X"96",X"84",X"74",X"6A",
		X"66",X"64",X"64",X"66",X"6A",X"6E",X"72",X"7A",X"84",X"8C",X"94",X"9A",X"9C",X"9E",X"9E",X"98",
		X"86",X"76",X"6C",X"66",X"64",X"64",X"66",X"6A",X"6C",X"70",X"78",X"82",X"8C",X"94",X"9A",X"9C",
		X"9E",X"9E",X"98",X"86",X"76",X"6C",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"78",X"84",X"8E",
		X"96",X"9A",X"9E",X"9E",X"9E",X"96",X"84",X"74",X"6A",X"66",X"64",X"64",X"66",X"6A",X"6E",X"72",
		X"7C",X"86",X"8E",X"96",X"9A",X"9E",X"9E",X"9E",X"94",X"80",X"72",X"6A",X"64",X"64",X"64",X"68",
		X"6A",X"6E",X"74",X"7E",X"88",X"90",X"96",X"9A",X"9E",X"9E",X"9C",X"8E",X"7C",X"6E",X"68",X"64",
		X"64",X"66",X"68",X"6C",X"70",X"76",X"82",X"8C",X"94",X"98",X"9C",X"9E",X"9E",X"98",X"88",X"76",
		X"6C",X"66",X"64",X"64",X"66",X"6A",X"6E",X"72",X"7C",X"86",X"90",X"96",X"9A",X"9E",X"9E",X"9C",
		X"90",X"7E",X"70",X"68",X"64",X"62",X"64",X"68",X"6C",X"70",X"78",X"82",X"8C",X"94",X"9A",X"9E",
		X"9E",X"9E",X"98",X"88",X"78",X"6C",X"66",X"64",X"64",X"66",X"6A",X"6E",X"72",X"7C",X"86",X"90",
		X"96",X"9A",X"9E",X"9E",X"9E",X"90",X"7C",X"70",X"68",X"64",X"64",X"64",X"68",X"6A",X"70",X"78",
		X"84",X"8C",X"94",X"9A",X"9C",X"9E",X"9E",X"96",X"84",X"74",X"6A",X"66",X"64",X"64",X"68",X"6A",
		X"6E",X"74",X"7E",X"8A",X"90",X"98",X"9C",X"9E",X"9E",X"9A",X"8A",X"7A",X"6E",X"66",X"64",X"64",
		X"66",X"68",X"6C",X"70",X"7C",X"86",X"90",X"96",X"9A",X"9E",X"9E",X"9C",X"90",X"7C",X"70",X"68",
		X"64",X"64",X"66",X"68",X"6C",X"70",X"78",X"84",X"8C",X"94",X"9A",X"9C",X"9E",X"9E",X"92",X"80",
		X"72",X"6A",X"64",X"64",X"64",X"68",X"6A",X"6E",X"76",X"82",X"8C",X"94",X"98",X"9C",X"9E",X"9E",
		X"96",X"82",X"74",X"6A",X"64",X"64",X"64",X"68",X"6A",X"6E",X"76",X"80",X"8A",X"92",X"98",X"9C",
		X"9E",X"9E",X"98",X"84",X"76",X"6C",X"66",X"64",X"64",X"66",X"6A",X"6E",X"76",X"80",X"8A",X"92",
		X"98",X"9C",X"9E",X"9E",X"98",X"86",X"76",X"6C",X"66",X"64",X"66",X"68",X"6A",X"6E",X"76",X"80",
		X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"98",X"86",X"76",X"6A",X"66",X"64",X"64",X"68",X"6A",X"6E",
		X"74",X"80",X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"98",X"86",X"76",X"6C",X"66",X"64",X"66",X"68",
		X"6C",X"6E",X"74",X"7C",X"88",X"90",X"96",X"9C",X"9E",X"9E",X"9C",X"90",X"7C",X"70",X"68",X"64",
		X"64",X"66",X"68",X"6C",X"70",X"74",X"7E",X"8A",X"92",X"98",X"9C",X"9E",X"A0",X"9C",X"8A",X"7A",
		X"6E",X"68",X"66",X"64",X"66",X"68",X"6C",X"70",X"74",X"7E",X"88",X"90",X"98",X"9C",X"9E",X"A0",
		X"9E",X"90",X"7E",X"72",X"68",X"66",X"64",X"66",X"68",X"6A",X"6E",X"72",X"78",X"80",X"8A",X"94",
		X"98",X"9C",X"9E",X"9E",X"9C",X"8E",X"7C",X"70",X"68",X"64",X"64",X"66",X"68",X"6C",X"6E",X"72",
		X"78",X"80",X"8A",X"94",X"98",X"9E",X"A0",X"A0",X"9E",X"90",X"7E",X"70",X"68",X"64",X"64",X"64",
		X"68",X"6A",X"6E",X"72",X"74",X"7C",X"86",X"90",X"96",X"9C",X"9E",X"A0",X"A0",X"9A",X"86",X"76",
		X"6C",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"72",X"78",X"7E",X"88",X"92",X"98",X"9C",X"A0",
		X"A0",X"A0",X"96",X"84",X"74",X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"78",X"7E",
		X"88",X"90",X"98",X"9C",X"A0",X"A0",X"A0",X"9A",X"88",X"76",X"6C",X"66",X"62",X"62",X"64",X"68",
		X"6C",X"70",X"72",X"76",X"7A",X"82",X"8C",X"94",X"9A",X"A0",X"A0",X"A0",X"A0",X"96",X"84",X"74",
		X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",X"6E",X"72",X"76",X"7A",X"82",X"8C",X"94",X"9A",X"9E",
		X"A0",X"A0",X"A0",X"96",X"82",X"74",X"6A",X"64",X"64",X"64",X"66",X"68",X"6C",X"70",X"72",X"76",
		X"7A",X"7E",X"88",X"90",X"98",X"9C",X"A0",X"A2",X"A2",X"9C",X"8C",X"7A",X"6E",X"66",X"64",X"62",
		X"64",X"68",X"6A",X"6E",X"70",X"74",X"78",X"7C",X"82",X"8C",X"94",X"9A",X"9E",X"A0",X"A0",X"A0",
		X"98",X"84",X"76",X"6C",X"66",X"64",X"62",X"64",X"68",X"6A",X"6E",X"72",X"74",X"78",X"7C",X"82",
		X"8C",X"94",X"9A",X"9E",X"A0",X"A0",X"A0",X"9A",X"8A",X"78",X"6C",X"66",X"64",X"62",X"64",X"66",
		X"6A",X"6C",X"70",X"74",X"76",X"7A",X"80",X"88",X"90",X"98",X"9E",X"A0",X"A2",X"A0",X"9E",X"90",
		X"7E",X"70",X"68",X"64",X"62",X"64",X"66",X"6A",X"6C",X"6E",X"72",X"76",X"78",X"7C",X"82",X"8A",
		X"94",X"9A",X"9E",X"A0",X"A2",X"A2",X"9C",X"8C",X"7A",X"6E",X"66",X"64",X"64",X"64",X"66",X"6A",
		X"6C",X"70",X"74",X"76",X"7A",X"7C",X"82",X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9C",X"8A",
		X"78",X"6C",X"66",X"64",X"62",X"64",X"66",X"6A",X"6C",X"70",X"74",X"76",X"7A",X"7E",X"82",X"8A",
		X"92",X"9A",X"9E",X"A2",X"A2",X"A2",X"9E",X"90",X"7E",X"70",X"68",X"64",X"62",X"64",X"64",X"68",
		X"6A",X"6E",X"72",X"76",X"7A",X"7C",X"7E",X"86",X"8E",X"96",X"9C",X"9E",X"A2",X"A2",X"A0",X"98",
		X"86",X"76",X"6C",X"66",X"62",X"62",X"64",X"66",X"6A",X"6C",X"70",X"74",X"78",X"7A",X"7E",X"80",
		X"88",X"92",X"98",X"9E",X"A0",X"A2",X"A2",X"A0",X"94",X"80",X"72",X"68",X"64",X"62",X"62",X"64",
		X"68",X"6A",X"6E",X"70",X"74",X"78",X"7A",X"7E",X"82",X"8A",X"92",X"98",X"9E",X"A0",X"A2",X"A2",
		X"9E",X"92",X"80",X"72",X"68",X"64",X"62",X"62",X"64",X"68",X"6A",X"6E",X"70",X"74",X"78",X"7A",
		X"7E",X"80",X"88",X"90",X"98",X"9E",X"A0",X"A2",X"A2",X"A0",X"96",X"84",X"74",X"6A",X"64",X"62",
		X"62",X"64",X"68",X"6A",X"6C",X"70",X"74",X"76",X"7A",X"7C",X"80",X"86",X"8E",X"96",X"9C",X"9E",
		X"A2",X"A2",X"A0",X"9A",X"88",X"78",X"6C",X"66",X"62",X"62",X"64",X"66",X"6A",X"6C",X"70",X"72",
		X"76",X"7A",X"7C",X"7E",X"82",X"8A",X"94",X"9A",X"9E",X"A0",X"A2",X"A2",X"9E",X"92",X"7E",X"70",
		X"66",X"62",X"60",X"62",X"64",X"66",X"6A",X"6E",X"72",X"74",X"78",X"7C",X"7E",X"80",X"86",X"8E",
		X"96",X"9C",X"A0",X"A2",X"A2",X"A0",X"9C",X"8C",X"7C",X"70",X"68",X"64",X"64",X"64",X"66",X"68",
		X"6C",X"6E",X"70",X"74",X"78",X"7A",X"7E",X"80",X"86",X"8E",X"96",X"9C",X"A0",X"A2",X"A2",X"A0",
		X"9C",X"8A",X"78",X"6C",X"66",X"62",X"62",X"64",X"66",X"68",X"6C",X"6E",X"72",X"76",X"78",X"7C",
		X"7E",X"80",X"86",X"90",X"96",X"9C",X"A0",X"A2",X"A2",X"A0",X"9A",X"8A",X"78",X"6C",X"66",X"64",
		X"62",X"64",X"66",X"68",X"6C",X"6E",X"72",X"74",X"78",X"7A",X"7E",X"80",X"84",X"8E",X"94",X"9A",
		X"A0",X"A2",X"A2",X"A2",X"9C",X"8C",X"7A",X"6E",X"66",X"62",X"62",X"62",X"64",X"68",X"6A",X"6E",
		X"70",X"74",X"76",X"7A",X"7E",X"80",X"84",X"8C",X"94",X"9A",X"9E",X"A0",X"A2",X"A0",X"9E",X"92",
		X"80",X"72",X"68",X"64",X"62",X"62",X"64",X"66",X"6A",X"6E",X"70",X"74",X"76",X"7A",X"7C",X"7E",
		X"82",X"88",X"90",X"98",X"9C",X"A0",X"A2",X"A2",X"A0",X"9A",X"88",X"76",X"6C",X"64",X"62",X"62",
		X"64",X"66",X"68",X"6C",X"6E",X"72",X"76",X"78",X"7C",X"7E",X"80",X"84",X"8C",X"94",X"9A",X"9E",
		X"A0",X"A2",X"A0",X"9E",X"90",X"7E",X"70",X"68",X"62",X"62",X"64",X"64",X"68",X"6C",X"6E",X"72",
		X"74",X"76",X"7A",X"7C",X"80",X"82",X"86",X"8E",X"96",X"9C",X"A0",X"A2",X"A2",X"A0",X"9C",X"8C",
		X"7A",X"6E",X"66",X"64",X"62",X"64",X"66",X"68",X"6C",X"6E",X"72",X"74",X"76",X"7A",X"7C",X"7E",
		X"82",X"88",X"90",X"98",X"9C",X"A0",X"A2",X"A0",X"A0",X"98",X"88",X"78",X"6C",X"66",X"62",X"62",
		X"64",X"66",X"68",X"6C",X"6E",X"72",X"76",X"78",X"7A",X"7E",X"82",X"88",X"92",X"98",X"9C",X"A0",
		X"A2",X"A0",X"9E",X"96",X"84",X"74",X"6A",X"64",X"62",X"62",X"64",X"66",X"68",X"6C",X"70",X"72",
		X"76",X"7A",X"7C",X"80",X"88",X"90",X"98",X"9C",X"A0",X"A2",X"A0",X"9E",X"96",X"84",X"74",X"6A",
		X"64",X"62",X"62",X"64",X"66",X"6A",X"6C",X"70",X"74",X"78",X"7A",X"7E",X"84",X"8C",X"94",X"9A",
		X"9E",X"A0",X"A0",X"9E",X"9A",X"88",X"78",X"6C",X"66",X"64",X"64",X"64",X"66",X"6A",X"6C",X"70",
		X"72",X"76",X"7A",X"7E",X"86",X"90",X"96",X"9C",X"9E",X"A0",X"A0",X"9E",X"96",X"84",X"74",X"6C",
		X"66",X"64",X"64",X"66",X"68",X"6A",X"6E",X"72",X"74",X"78",X"7C",X"82",X"8C",X"94",X"9A",X"9E",
		X"A0",X"A0",X"A0",X"98",X"86",X"76",X"6C",X"66",X"62",X"62",X"64",X"68",X"6A",X"6E",X"72",X"76",
		X"78",X"7E",X"86",X"90",X"98",X"9C",X"A0",X"A0",X"A0",X"9C",X"92",X"80",X"72",X"6A",X"66",X"64",
		X"64",X"66",X"6A",X"6C",X"70",X"74",X"78",X"7A",X"82",X"8C",X"94",X"9A",X"9E",X"A0",X"9E",X"9C",
		X"94",X"82",X"74",X"6A",X"66",X"64",X"64",X"66",X"68",X"6C",X"70",X"74",X"76",X"7C",X"84",X"8E",
		X"96",X"9C",X"9E",X"A0",X"9E",X"9C",X"90",X"7E",X"72",X"68",X"66",X"64",X"64",X"68",X"6A",X"6E",
		X"70",X"74",X"78",X"7E",X"88",X"92",X"98",X"9C",X"9E",X"A0",X"9E",X"98",X"88",X"78",X"6C",X"66",
		X"64",X"64",X"66",X"68",X"6A",X"6E",X"72",X"76",X"7C",X"86",X"90",X"96",X"9A",X"9E",X"9E",X"9C",
		X"98",X"8A",X"7A",X"6E",X"68",X"64",X"64",X"66",X"68",X"6A",X"6E",X"72",X"76",X"7C",X"86",X"90",
		X"96",X"9C",X"9E",X"9E",X"9E",X"98",X"88",X"78",X"6E",X"68",X"64",X"64",X"66",X"6A",X"6C",X"70",
		X"74",X"78",X"80",X"8A",X"92",X"98",X"9C",X"9E",X"9E",X"9C",X"92",X"80",X"74",X"6C",X"66",X"66",
		X"66",X"68",X"6A",X"6E",X"72",X"74",X"7A",X"86",X"8E",X"94",X"9A",X"9C",X"9C",X"9A",X"96",X"88",
		X"78",X"6E",X"68",X"66",X"66",X"68",X"6A",X"6C",X"70",X"74",X"78",X"82",X"8C",X"94",X"9A",X"9C",
		X"9E",X"9C",X"98",X"8C",X"7A",X"70",X"6A",X"66",X"64",X"66",X"6A",X"6C",X"70",X"74",X"78",X"82",
		X"8C",X"94",X"9A",X"9C",X"9E",X"9C",X"98",X"8A",X"7C",X"70",X"6A",X"66",X"66",X"66",X"68",X"6C",
		X"70",X"74",X"7A",X"84",X"8C",X"94",X"9A",X"9C",X"9E",X"9C",X"96",X"88",X"78",X"6E",X"68",X"66",
		X"66",X"68",X"6A",X"6E",X"70",X"74",X"7C",X"86",X"90",X"96",X"9A",X"9C",X"9C",X"9A",X"92",X"82",
		X"74",X"6C",X"68",X"66",X"66",X"68",X"6C",X"6E",X"72",X"78",X"82",X"8C",X"94",X"98",X"9C",X"9C",
		X"9C",X"96",X"8A",X"7A",X"70",X"6A",X"66",X"66",X"68",X"6A",X"6E",X"70",X"74",X"7C",X"88",X"90",
		X"96",X"9A",X"9C",X"9C",X"98",X"90",X"7E",X"72",X"6A",X"66",X"66",X"66",X"6A",X"6C",X"70",X"74",
		X"7A",X"84",X"8E",X"94",X"98",X"9C",X"9C",X"9A",X"92",X"84",X"76",X"6C",X"68",X"66",X"66",X"68",
		X"6C",X"6E",X"72",X"78",X"82",X"8C",X"94",X"98",X"9A",X"9C",X"9A",X"94",X"86",X"78",X"6E",X"68",
		X"68",X"68",X"6A",X"6C",X"6E",X"72",X"78",X"82",X"8C",X"94",X"98",X"9A",X"9A",X"9A",X"94",X"86",
		X"78",X"6E",X"68",X"66",X"66",X"68",X"6C",X"6E",X"72",X"7A",X"84",X"8C",X"94",X"98",X"9A",X"9A",
		X"98",X"92",X"82",X"76",X"6C",X"68",X"68",X"68",X"6A",X"6E",X"70",X"74",X"7C",X"86",X"8E",X"96",
		X"9A",X"9C",X"9A",X"98",X"90",X"80",X"74",X"6C",X"68",X"66",X"66",X"6A",X"6C",X"70",X"74",X"7E",
		X"88",X"90",X"96",X"9A",X"9A",X"98",X"96",X"8C",X"7C",X"72",X"6A",X"68",X"68",X"68",X"6A",X"6E",
		X"70",X"76",X"80",X"8A",X"92",X"98",X"9A",X"9A",X"98",X"94",X"88",X"78",X"70",X"6A",X"68",X"68",
		X"68",X"6C",X"70",X"72",X"7A",X"84",X"8E",X"94",X"98",X"9A",X"9A",X"96",X"90",X"82",X"74",X"6E",
		X"68",X"68",X"68",X"6A",X"6C",X"70",X"74",X"7E",X"88",X"90",X"96",X"9A",X"9A",X"98",X"94",X"8A",
		X"7A",X"70",X"6A",X"68",X"66",X"6A",X"6C",X"6E",X"72",X"7A",X"84",X"8C",X"94",X"98",X"9A",X"98",
		X"96",X"8E",X"80",X"74",X"6C",X"68",X"68",X"68",X"6A",X"6E",X"70",X"76",X"80",X"8A",X"92",X"96",
		X"9A",X"9A",X"98",X"92",X"84",X"76",X"6E",X"68",X"68",X"68",X"6A",X"6C",X"70",X"74",X"7E",X"88",
		X"90",X"96",X"98",X"9A",X"98",X"94",X"8A",X"7A",X"70",X"6A",X"68",X"68",X"68",X"6C",X"6E",X"72",
		X"7A",X"86",X"8E",X"94",X"98",X"9A",X"98",X"96",X"8C",X"7E",X"72",X"6C",X"68",X"68",X"6A",X"6C",
		X"6E",X"70",X"78",X"84",X"8C",X"92",X"96",X"98",X"98",X"96",X"90",X"80",X"74",X"6E",X"6A",X"68",
		X"6A",X"6C",X"6E",X"72",X"78",X"82",X"8C",X"92",X"96",X"98",X"98",X"96",X"90",X"82",X"76",X"6E",
		X"6A",X"68",X"6A",X"6C",X"6E",X"70",X"76",X"80",X"8A",X"92",X"96",X"98",X"98",X"96",X"90",X"82",
		X"76",X"6E",X"6A",X"68",X"6A",X"6C",X"6E",X"72",X"78",X"82",X"8C",X"92",X"96",X"98",X"98",X"96",
		X"90",X"80",X"76",X"6E",X"6A",X"6A",X"6A",X"6C",X"6E",X"72",X"78",X"82",X"8A",X"92",X"96",X"98",
		X"98",X"96",X"90",X"82",X"76",X"6E",X"6A",X"6A",X"6A",X"6C",X"6E",X"72",X"76",X"82",X"8C",X"92",
		X"96",X"98",X"96",X"94",X"8C",X"7E",X"74",X"6C",X"6A",X"6A",X"6A",X"6C",X"6E",X"72",X"78",X"80",
		X"8A",X"92",X"96",X"98",X"98",X"96",X"90",X"84",X"76",X"6E",X"6A",X"6A",X"6A",X"6C",X"6E",X"70",
		X"74",X"7A",X"84",X"8C",X"94",X"98",X"9A",X"98",X"96",X"90",X"82",X"76",X"6E",X"6A",X"6A",X"6A",
		X"6C",X"6E",X"72",X"74",X"78",X"82",X"8C",X"92",X"96",X"98",X"98",X"96",X"90",X"84",X"78",X"70",
		X"6C",X"6A",X"6A",X"6C",X"6E",X"70",X"74",X"76",X"7E",X"88",X"90",X"94",X"98",X"98",X"96",X"94",
		X"8C",X"7E",X"74",X"6C",X"6A",X"68",X"6A",X"6C",X"6E",X"70",X"74",X"78",X"7E",X"88",X"92",X"98",
		X"9A",X"9A",X"98",X"96",X"8C",X"80",X"74",X"6E",X"6C",X"6A",X"6A",X"6C",X"6E",X"72",X"74",X"78",
		X"7C",X"86",X"8E",X"94",X"98",X"9A",X"98",X"96",X"90",X"84",X"78",X"70",X"6C",X"6A",X"6A",X"6A",
		X"6C",X"6E",X"72",X"74",X"78",X"7C",X"86",X"8E",X"96",X"98",X"9A",X"98",X"96",X"90",X"84",X"76",
		X"70",X"6A",X"6A",X"6A",X"6C",X"6E",X"70",X"72",X"76",X"78",X"7C",X"86",X"8E",X"94",X"98",X"9A",
		X"98",X"96",X"90",X"86",X"7A",X"72",X"6C",X"6A",X"6A",X"6C",X"6E",X"70",X"72",X"74",X"78",X"7A",
		X"80",X"8A",X"90",X"96",X"9A",X"9A",X"98",X"94",X"8E",X"82",X"76",X"70",X"6C",X"6A",X"6A",X"6C",
		X"6E",X"70",X"72",X"76",X"78",X"7A",X"80",X"8A",X"92",X"96",X"9A",X"98",X"98",X"94",X"8E",X"80",
		X"76",X"6E",X"6A",X"6A",X"6A",X"6C",X"6E",X"70",X"72",X"76",X"78",X"7A",X"7E",X"88",X"90",X"96",
		X"98",X"9A",X"98",X"96",X"90",X"86",X"7A",X"70",X"6C",X"6A",X"68",X"6A",X"6C",X"6E",X"72",X"74",
		X"78",X"7A",X"7C",X"82",X"8C",X"92",X"96",X"9A",X"9A",X"96",X"94",X"8E",X"82",X"76",X"70",X"6C",
		X"6A",X"6A",X"6C",X"6E",X"70",X"72",X"74",X"76",X"7A",X"7C",X"80",X"8A",X"92",X"96",X"98",X"98",
		X"98",X"94",X"90",X"84",X"78",X"72",X"6C",X"6C",X"6A",X"6C",X"6E",X"70",X"72",X"76",X"78",X"7A",
		X"7C",X"80",X"88",X"90",X"96",X"98",X"98",X"98",X"96",X"92",X"88",X"7C",X"72",X"6E",X"6C",X"6A",
		X"6C",X"6C",X"6E",X"72",X"74",X"76",X"78",X"7C",X"7E",X"82",X"8A",X"92",X"96",X"98",X"98",X"96",
		X"94",X"8E",X"84",X"78",X"72",X"6C",X"6C",X"6A",X"6C",X"6E",X"70",X"72",X"74",X"76",X"7A",X"7C",
		X"7E",X"82",X"8C",X"92",X"96",X"9A",X"98",X"96",X"94",X"8E",X"84",X"78",X"70",X"6C",X"6A",X"6A",
		X"6C",X"6E",X"70",X"72",X"74",X"76",X"7A",X"7C",X"7E",X"82",X"8A",X"92",X"96",X"98",X"98",X"96",
		X"94",X"90",X"86",X"7A",X"72",X"6E",X"6C",X"6A",X"6C",X"6C",X"6E",X"72",X"74",X"76",X"78",X"7C",
		X"7E",X"80",X"86",X"8E",X"94",X"98",X"98",X"98",X"94",X"92",X"8A",X"7E",X"74",X"6E",X"6C",X"6A",
		X"6C",X"6C",X"6E",X"70",X"72",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"88",X"90",X"94",X"98",X"98",
		X"96",X"94",X"90",X"88",X"7C",X"74",X"6E",X"6C",X"6C",X"6C",X"6E",X"70",X"72",X"74",X"76",X"78",
		X"7A",X"7C",X"7E",X"82",X"8A",X"90",X"96",X"98",X"98",X"96",X"92",X"8E",X"86",X"7A",X"72",X"6E",
		X"6A",X"6A",X"6C",X"6C",X"6E",X"72",X"74",X"76",X"7A",X"7C",X"7E",X"80",X"82",X"88",X"90",X"94",
		X"98",X"98",X"96",X"94",X"90",X"88",X"7E",X"74",X"70",X"6E",X"6C",X"6C",X"6E",X"70",X"72",X"74",
		X"76",X"78",X"7A",X"7C",X"7E",X"80",X"84",X"8C",X"92",X"96",X"96",X"96",X"94",X"90",X"8C",X"82",
		X"78",X"70",X"6E",X"6C",X"6C",X"6E",X"6E",X"70",X"72",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"80",
		X"88",X"90",X"94",X"96",X"96",X"96",X"94",X"90",X"88",X"7E",X"74",X"70",X"6C",X"6C",X"6C",X"6E",
		X"70",X"72",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"84",X"8A",X"90",X"96",X"96",X"96",X"94",
		X"92",X"8E",X"84",X"7A",X"74",X"70",X"6E",X"6C",X"6C",X"6E",X"70",X"72",X"74",X"76",X"78",X"7A",
		X"7C",X"7E",X"80",X"84",X"8C",X"92",X"96",X"96",X"94",X"94",X"90",X"8C",X"82",X"78",X"72",X"6E",
		X"6E",X"6C",X"6E",X"70",X"70",X"72",X"74",X"78",X"78",X"7C",X"7C",X"7E",X"80",X"84",X"8C",X"92",
		X"96",X"96",X"96",X"94",X"90",X"8C",X"82",X"78",X"72",X"6E",X"6E",X"6E",X"6E",X"70",X"70",X"72",
		X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"84",X"8A",X"92",X"94",X"96",X"96",X"94",X"90",X"8C",
		X"84",X"7A",X"72",X"6E",X"6C",X"6C",X"6E",X"6E",X"70",X"72",X"74",X"78",X"7A",X"7C",X"7E",X"7E",
		X"80",X"84",X"8A",X"90",X"94",X"96",X"96",X"94",X"90",X"8E",X"86",X"7C",X"76",X"70",X"6E",X"6E",
		X"6E",X"70",X"72",X"72",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"86",X"8E",X"92",X"94",
		X"94",X"94",X"90",X"8E",X"8A",X"80",X"78",X"72",X"70",X"6E",X"6E",X"70",X"70",X"72",X"74",X"76",
		X"78",X"7A",X"7C",X"7E",X"80",X"80",X"82",X"88",X"8E",X"92",X"94",X"94",X"92",X"90",X"8C",X"86",
		X"7C",X"76",X"72",X"6E",X"6E",X"6E",X"70",X"72",X"72",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",
		X"80",X"84",X"8C",X"90",X"94",X"94",X"94",X"92",X"8E",X"8A",X"82",X"7A",X"74",X"70",X"6E",X"6E",
		X"6E",X"70",X"72",X"74",X"76",X"78",X"7A",X"7C",X"7C",X"7E",X"80",X"82",X"86",X"8C",X"92",X"94",
		X"94",X"92",X"90",X"8E",X"88",X"80",X"78",X"72",X"70",X"6E",X"6E",X"70",X"70",X"72",X"74",X"76",
		X"78",X"7A",X"7C",X"7E",X"7E",X"80",X"86",X"8C",X"90",X"94",X"92",X"92",X"90",X"8C",X"88",X"7E",
		X"78",X"72",X"70",X"70",X"6E",X"70",X"72",X"72",X"74",X"78",X"78",X"7A",X"7C",X"7E",X"80",X"86",
		X"8C",X"90",X"92",X"92",X"92",X"8E",X"8C",X"86",X"7E",X"76",X"72",X"6E",X"6E",X"70",X"70",X"72",
		X"74",X"76",X"78",X"7A",X"7C",X"7E",X"80",X"82",X"8A",X"90",X"92",X"92",X"92",X"90",X"8C",X"8A",
		X"82",X"7A",X"74",X"72",X"70",X"70",X"70",X"72",X"74",X"76",X"78",X"7A",X"7A",X"7C",X"7E",X"84",
		X"8A",X"90",X"92",X"92",X"90",X"8E",X"8C",X"88",X"80",X"78",X"74",X"72",X"70",X"70",X"72",X"72",
		X"74",X"76",X"78",X"7A",X"7A",X"7E",X"82",X"88",X"8E",X"90",X"92",X"90",X"8E",X"8C",X"88",X"82",
		X"7A",X"74",X"72",X"70",X"70",X"72",X"72",X"74",X"76",X"78",X"7A",X"7C",X"7E",X"82",X"8A",X"8E",
		X"90",X"90",X"90",X"8E",X"8A",X"86",X"7E",X"78",X"74",X"72",X"70",X"72",X"72",X"74",X"76",X"78",
		X"7A",X"7C",X"7C",X"80",X"88",X"8C",X"90",X"90",X"8E",X"8E",X"8C",X"88",X"80",X"7A",X"74",X"72",
		X"70",X"70",X"72",X"74",X"76",X"76",X"78",X"7A",X"7C",X"82",X"88",X"8C",X"90",X"90",X"8E",X"8C",
		X"8A",X"86",X"80",X"78",X"74",X"72",X"70",X"72",X"72",X"74",X"74",X"76",X"7A",X"7A",X"7E",X"84",
		X"8A",X"8E",X"90",X"90",X"8E",X"8C",X"88",X"82",X"7C",X"76",X"74",X"72",X"72",X"72",X"74",X"76",
		X"76",X"78",X"7A",X"7C",X"82",X"88",X"8E",X"8E",X"8E",X"8E",X"8C",X"8A",X"84",X"7C",X"76",X"72",
		X"72",X"72",X"72",X"74",X"76",X"78",X"7A",X"7A",X"7C",X"84",X"88",X"8C",X"8E",X"8E",X"8E",X"8A",
		X"8A",X"84",X"7C",X"78",X"74",X"72",X"72",X"72",X"74",X"76",X"76",X"7A",X"7A",X"7E",X"84",X"8A",
		X"8C",X"8E",X"8C",X"8C",X"8A",X"86",X"80",X"7A",X"76",X"74",X"72",X"74",X"74",X"76",X"76",X"78",
		X"7A",X"7C",X"80",X"88",X"8C",X"8E",X"8E",X"8C",X"8A",X"88",X"84",X"7C",X"78",X"74",X"74",X"72",
		X"74",X"74",X"76",X"78",X"7A",X"7C",X"80",X"86",X"8A",X"8C",X"8E",X"8C",X"8C",X"88",X"86",X"80",
		X"78",X"76",X"74",X"72",X"72",X"74",X"76",X"76",X"78",X"7A",X"7E",X"86",X"8A",X"8C",X"8C",X"8C",
		X"8A",X"88",X"86",X"80",X"7A",X"76",X"74",X"74",X"74",X"74",X"76",X"78",X"7A",X"7C",X"80",X"86",
		X"8A",X"8C",X"8C",X"8C",X"8A",X"88",X"84",X"7E",X"7A",X"76",X"74",X"74",X"74",X"74",X"76",X"78",
		X"7A",X"7A",X"80",X"86",X"8A",X"8C",X"8C",X"8C",X"8A",X"88",X"82",X"7C",X"78",X"74",X"74",X"74",
		X"74",X"76",X"76",X"78",X"7A",X"7E",X"84",X"88",X"8A",X"8C",X"8C",X"8A",X"88",X"86",X"80",X"7A",
		X"76",X"74",X"74",X"74",X"76",X"76",X"78",X"7A",X"7C",X"82",X"86",X"8A",X"8A",X"8A",X"8A",X"88",
		X"86",X"80",X"7A",X"76",X"76",X"74",X"74",X"76",X"76",X"78",X"78",X"7A",X"80",X"86",X"8A",X"8C",
		X"8C",X"8A",X"88",X"86",X"82",X"7C",X"78",X"76",X"74",X"74",X"76",X"76",X"78",X"78",X"7A",X"80",
		X"86",X"88",X"8A",X"8C",X"8A",X"8A",X"86",X"84",X"7E",X"78",X"76",X"74",X"74",X"76",X"76",X"78",
		X"7A",X"7A",X"7E",X"84",X"88",X"8A",X"8A",X"8A",X"8A",X"88",X"84",X"7E",X"78",X"76",X"74",X"76",
		X"76",X"76",X"78",X"7A",X"7C",X"80",X"86",X"88",X"8A",X"8A",X"8A",X"88",X"86",X"82",X"7C",X"78",
		X"76",X"76",X"74",X"76",X"78",X"78",X"7A",X"7C",X"82",X"86",X"88",X"8A",X"8A",X"88",X"88",X"84",
		X"82",X"7C",X"78",X"76",X"76",X"76",X"76",X"78",X"78",X"7A",X"7C",X"82",X"86",X"88",X"8A",X"8A",
		X"88",X"86",X"84",X"80",X"7A",X"78",X"76",X"76",X"76",X"76",X"78",X"7A",X"7A",X"7E",X"84",X"88",
		X"8A",X"88",X"88",X"88",X"86",X"82",X"7E",X"7A",X"76",X"76",X"76",X"76",X"78",X"78",X"7A",X"7C",
		X"82",X"86",X"88",X"8A",X"8A",X"88",X"86",X"84",X"80",X"7C",X"78",X"76",X"76",X"76",X"76",X"78",
		X"7A",X"7A",X"7E",X"84",X"86",X"88",X"8A",X"88",X"86",X"86",X"82",X"7E",X"7A",X"76",X"76",X"76",
		X"76",X"78",X"78",X"78",X"7C",X"82",X"86",X"88",X"8A",X"88",X"88",X"86",X"84",X"80",X"7C",X"78",
		X"76",X"76",X"78",X"78",X"78",X"7A",X"7C",X"80",X"84",X"88",X"88",X"88",X"88",X"86",X"84",X"82",
		X"7C",X"78",X"76",X"76",X"76",X"78",X"78",X"7A",X"7C",X"80",X"84",X"86",X"88",X"88",X"88",X"86",
		X"84",X"80",X"7C",X"7A",X"76",X"76",X"76",X"76",X"78",X"7A",X"7A",X"7E",X"84",X"86",X"88",X"88",
		X"88",X"86",X"84",X"82",X"7E",X"7A",X"78",X"76",X"76",X"78",X"78",X"7A",X"7A",X"7E",X"84",X"86",
		X"88",X"88",X"88",X"88",X"86",X"82",X"7E",X"7A",X"78",X"78",X"76",X"78",X"78",X"7A",X"7A",X"7E",
		X"82",X"86",X"88",X"88",X"88",X"86",X"86",X"82",X"7E",X"7C",X"78",X"78",X"78",X"76",X"78",X"7A",
		X"7A",X"7E",X"82",X"86",X"86",X"88",X"88",X"86",X"86",X"82",X"7E",X"7A",X"78",X"78",X"78",X"78",
		X"78",X"7A",X"7A",X"7C",X"82",X"84",X"86",X"88",X"86",X"86",X"84",X"82",X"7E",X"7A",X"78",X"78",
		X"78",X"78",X"78",X"78",X"7A",X"7E",X"82",X"86",X"88",X"88",X"88",X"86",X"86",X"82",X"7E",X"7C",
		X"7A",X"78",X"78",X"78",X"78",X"7A",X"7A",X"7E",X"82",X"84",X"86",X"86",X"86",X"86",X"84",X"82",
		X"7E",X"7A",X"78",X"76",X"76",X"76",X"78",X"78",X"7A",X"7C",X"82",X"86",X"88",X"88",X"88",X"88",
		X"86",X"84",X"80",X"7C",X"7A",X"78",X"78",X"78",X"7A",X"7A",X"7A",X"7C",X"7E",X"82",X"86",X"86",
		X"88",X"88",X"86",X"84",X"82",X"7E",X"7A",X"78",X"78",X"78",X"78",X"78",X"7A",X"7A",X"7C",X"7E",
		X"82",X"84",X"86",X"86",X"86",X"86",X"84",X"82",X"7E",X"7C",X"7A",X"78",X"78",X"78",X"7A",X"7A",
		X"7A",X"7C",X"7E",X"80",X"84",X"86",X"88",X"88",X"86",X"86",X"84",X"82",X"7E",X"7A",X"7A",X"78",
		X"78",X"78",X"7A",X"7A",X"7A",X"7C",X"7C",X"80",X"84",X"86",X"88",X"88",X"86",X"84",X"84",X"82",
		X"7E",X"7C",X"7A",X"78",X"78",X"78",X"7A",X"7A",X"7A",X"7C",X"7C",X"7E",X"82",X"84",X"86",X"86",
		X"86",X"86",X"84",X"82",X"80",X"7C",X"7A",X"7A",X"78",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",X"7C",
		X"7E",X"82",X"84",X"86",X"88",X"86",X"86",X"86",X"84",X"80",X"7C",X"7A",X"78",X"78",X"78",X"7A",
		X"7A",X"7A",X"7C",X"7C",X"7C",X"7E",X"82",X"84",X"86",X"86",X"86",X"86",X"84",X"82",X"80",X"7C",
		X"7A",X"7A",X"78",X"78",X"7A",X"7A",X"7A",X"7A",X"7C",X"7E",X"7E",X"80",X"82",X"86",X"86",X"86",
		X"86",X"86",X"84",X"82",X"7E",X"7C",X"7A",X"78",X"78",X"78",X"78",X"78",X"7A",X"7A",X"7C",X"7E",
		X"7E",X"80",X"84",X"86",X"88",X"88",X"88",X"86",X"84",X"82",X"80",X"7C",X"7A",X"7A",X"7A",X"7A",
		X"7A",X"7A",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"82",X"84",X"86",X"86",X"86",X"84",X"84",X"82",
		X"80",X"7E",X"7A",X"78",X"78",X"78",X"7A",X"7A",X"7A",X"7C",X"7C",X"7E",X"7E",X"7E",X"80",X"84",
		X"86",X"86",X"86",X"86",X"84",X"84",X"82",X"80",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",
		X"7C",X"7C",X"7E",X"7E",X"7E",X"80",X"84",X"86",X"86",X"86",X"86",X"84",X"84",X"82",X"80",X"7C",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"80",X"82",X"84",X"86",
		X"86",X"86",X"84",X"84",X"82",X"80",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",
		X"7C",X"7E",X"7E",X"7E",X"80",X"82",X"86",X"86",X"86",X"86",X"84",X"84",X"82",X"7E",X"7C",X"7A",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"80",X"84",X"84",X"86",
		X"86",X"84",X"84",X"82",X"82",X"7E",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",
		X"7E",X"7E",X"7E",X"80",X"82",X"84",X"86",X"86",X"84",X"84",X"82",X"82",X"82",X"7E",X"7C",X"7A",
		X"7A",X"78",X"7A",X"7A",X"7A",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"82",X"84",X"84",
		X"84",X"84",X"84",X"82",X"82",X"80",X"7E",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",
		X"7E",X"7E",X"7E",X"80",X"80",X"80",X"82",X"84",X"84",X"84",X"84",X"82",X"82",X"82",X"7E",X"7C",
		X"7C",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"80",X"7E",X"7E",X"82",X"84",
		X"84",X"84",X"84",X"84",X"84",X"82",X"80",X"7E",X"7C",X"7C",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"82",X"84",X"84",X"84",X"84",X"84",X"84",X"82",X"80",
		X"7E",X"7C",X"7C",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",
		X"80",X"82",X"84",X"84",X"84",X"84",X"82",X"82",X"80",X"7E",X"7C",X"7C",X"7C",X"7A",X"7A",X"7A",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"80",X"82",X"84",X"84",X"84",X"84",X"84",
		X"82",X"82",X"80",X"7E",X"7C",X"7C",X"7C",X"7A",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"80",X"80",X"82",X"84",X"84",X"84",X"84",X"82",X"82",X"80",X"7E",X"7C",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"82",X"84",X"84",
		X"84",X"84",X"84",X"82",X"82",X"80",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"82",X"82",X"84",X"82",X"82",X"82",X"82",X"80",
		X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",
		X"80",X"80",X"82",X"82",X"84",X"82",X"82",X"82",X"82",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"7E",X"80",X"80",X"82",X"82",X"84",X"84",
		X"82",X"82",X"82",X"80",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"80",X"7E",X"80",X"80",X"82",X"84",X"84",X"84",X"82",X"82",X"80",X"80",X"7E",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",
		X"80",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"7E",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"82",X"82",X"84",X"84",X"82",
		X"82",X"82",X"80",X"80",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"7E",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"80",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"80",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7E",X"7C",X"7E",X"7E",X"7E",X"80",X"7E",X"80",X"80",X"80",X"82",X"82",X"82",X"82",X"82",X"80",
		X"80",X"80",X"7E",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"80",X"80",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"7E",X"7E",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"82",X"82",X"82",X"82",X"82",
		X"80",X"80",X"7E",X"7E",X"7E",X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",
		X"80",X"80",X"82",X"82",X"82",X"82",X"80",X"80",X"80",X"7E",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"82",X"82",X"82",X"82",X"80",X"80",X"80",
		X"7E",X"7E",X"7C",X"7C",X"7C",X"7C",X"7C",X"7E",X"7E",X"7C",X"7E",X"7E",X"7E",X"80",X"80",X"82",
		X"82",X"82",X"82",X"82",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"80",X"80",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"7E",X"7E",X"7E",X"7C",
		X"7C",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"82",X"82",X"82",X"82",X"82",
		X"80",X"7E",X"7E",X"7E",X"7E",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"82",
		X"82",X"82",X"82",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7C",X"7C",X"7E",X"7C",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"80",X"80",X"80",X"82",X"82",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7C",X"7E",
		X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"82",X"82",X"82",X"80",X"80",X"80",
		X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",
		X"82",X"82",X"82",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"80",X"80",X"80",X"82",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7C",X"7C",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"82",X"82",X"80",X"80",X"80",X"80",X"80",X"7E",X"7C",X"7C",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"80",X"80",X"80",X"82",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",
		X"82",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7C",X"7E",X"7E",
		X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7C",X"7C",X"7E",X"7C",
		X"7C",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"82",X"82",X"82",X"82",X"80",X"80",X"80",X"7E",X"7C",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",
		X"7E",X"7E",X"7C",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7E",X"7E",X"7C",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"82",X"80",X"80",
		X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7E",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7E",X"7E",X"7E",X"7E",X"7E",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"80",X"80",X"7F",X"7F",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"80",X"7F",X"80",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"7F",
		X"7F",X"7F",X"7F",X"80",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"80",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"83",X"83",X"84",X"84",X"84",
		X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"83",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",
		X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"79",X"77",X"76",X"74",X"73",X"73",X"74",X"74",X"76",X"77",
		X"77",X"7A",X"7A",X"7D",X"7F",X"80",X"81",X"81",X"83",X"84",X"86",X"87",X"87",X"87",X"89",X"89",
		X"89",X"89",X"89",X"87",X"87",X"87",X"87",X"87",X"86",X"86",X"86",X"84",X"84",X"84",X"83",X"83",
		X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"83",X"87",X"8A",X"8C",X"8D",X"8D",X"8C",X"8A",
		X"87",X"84",X"83",X"80",X"7D",X"7A",X"77",X"74",X"73",X"71",X"70",X"6E",X"6D",X"6D",X"6B",X"6B",
		X"6B",X"6B",X"6D",X"6D",X"6D",X"6E",X"70",X"70",X"70",X"6E",X"6B",X"6A",X"68",X"68",X"68",X"6A",
		X"6B",X"6E",X"71",X"74",X"77",X"7A",X"7F",X"81",X"84",X"89",X"8A",X"8D",X"90",X"93",X"95",X"96",
		X"98",X"99",X"9B",X"9B",X"9B",X"9B",X"99",X"99",X"99",X"98",X"96",X"96",X"95",X"93",X"92",X"93",
		X"96",X"9B",X"9F",X"A1",X"A1",X"A1",X"9E",X"99",X"95",X"8F",X"89",X"84",X"7F",X"79",X"73",X"6E",
		X"6A",X"67",X"62",X"61",X"5E",X"5C",X"5B",X"59",X"59",X"59",X"59",X"5B",X"5B",X"5C",X"5E",X"5F",
		X"62",X"64",X"67",X"68",X"6B",X"6E",X"70",X"73",X"76",X"77",X"7A",X"7C",X"7D",X"80",X"81",X"83",
		X"84",X"86",X"87",X"89",X"89",X"8A",X"8A",X"8C",X"8C",X"8D",X"8D",X"8D",X"8D",X"8D",X"8D",X"8C",
		X"8C",X"8C",X"89",X"84",X"81",X"7D",X"7A",X"79",X"79",X"77",X"79",X"79",X"7A",X"7C",X"7D",X"7F",
		X"80",X"81",X"84",X"86",X"87",X"89",X"8A",X"8A",X"8C",X"8D",X"8D",X"8F",X"8F",X"8F",X"8F",X"8F",
		X"8F",X"8F",X"8F",X"8D",X"8D",X"8D",X"8C",X"8A",X"8A",X"89",X"89",X"87",X"87",X"87",X"86",X"86",
		X"86",X"87",X"8F",X"96",X"9C",X"A2",X"A4",X"A4",X"9F",X"9B",X"96",X"8F",X"89",X"81",X"7A",X"74",
		X"6E",X"68",X"62",X"5E",X"59",X"56",X"55",X"52",X"50",X"50",X"50",X"50",X"50",X"52",X"53",X"55",
		X"56",X"59",X"5B",X"59",X"58",X"58",X"58",X"59",X"5C",X"5F",X"62",X"67",X"6B",X"70",X"74",X"79",
		X"7F",X"83",X"87",X"8A",X"8F",X"92",X"96",X"99",X"9C",X"9E",X"A1",X"A2",X"A4",X"A5",X"AA",X"B3",
		X"BA",X"C0",X"C3",X"C5",X"C3",X"C0",X"BC",X"B6",X"B0",X"A8",X"A1",X"99",X"92",X"8A",X"84",X"7D",
		X"79",X"73",X"6E",X"6A",X"67",X"64",X"61",X"5F",X"5E",X"5C",X"5C",X"5C",X"5C",X"5C",X"5E",X"5F",
		X"5F",X"61",X"62",X"64",X"67",X"68",X"6A",X"6D",X"6E",X"71",X"73",X"76",X"77",X"79",X"7A",X"7C",
		X"7D",X"7F",X"80",X"7D",X"7A",X"79",X"77",X"77",X"77",X"77",X"79",X"7A",X"7C",X"7F",X"80",X"83",
		X"86",X"87",X"8A",X"8C",X"8F",X"90",X"92",X"93",X"95",X"95",X"96",X"96",X"98",X"98",X"98",X"99",
		X"99",X"9E",X"A4",X"AA",X"B0",X"B3",X"B3",X"B1",X"AE",X"AA",X"A4",X"9E",X"96",X"90",X"89",X"83",
		X"7C",X"76",X"71",X"6B",X"67",X"64",X"61",X"5E",X"5B",X"59",X"58",X"58",X"58",X"58",X"58",X"58",
		X"59",X"5B",X"5C",X"5E",X"5F",X"5F",X"5E",X"5C",X"5C",X"5C",X"5E",X"61",X"62",X"65",X"6A",X"6D",
		X"71",X"74",X"79",X"7D",X"81",X"84",X"87",X"8C",X"8F",X"92",X"93",X"96",X"98",X"99",X"9B",X"9B",
		X"9C",X"9C",X"9C",X"9C",X"9C",X"9C",X"9B",X"99",X"99",X"98",X"96",X"95",X"95",X"93",X"92",X"90",
		X"90",X"95",X"9B",X"A2",X"A7",X"AA",X"AB",X"A8",X"A5",X"9F",X"98",X"92",X"8A",X"81",X"7C",X"74",
		X"6E",X"68",X"62",X"5E",X"5B",X"56",X"55",X"53",X"52",X"50",X"50",X"50",X"50",X"52",X"53",X"55",
		X"56",X"59",X"5B",X"5E",X"61",X"64",X"67",X"6A",X"6D",X"70",X"73",X"76",X"79",X"7C",X"7D",X"80",
		X"83",X"84",X"86",X"89",X"8A",X"8C",X"8C",X"8D",X"8F",X"90",X"90",X"92",X"92",X"92",X"92",X"92",
		X"90",X"90",X"8F",X"8D",X"89",X"84",X"81",X"7F",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7F",
		X"80",X"81",X"84",X"86",X"87",X"89",X"8A",X"8C",X"8D",X"8D",X"8F",X"8F",X"90",X"90",X"90",X"90",
		X"90",X"90",X"8F",X"8F",X"8D",X"8D",X"8C",X"8C",X"8A",X"8A",X"89",X"87",X"86",X"84",X"84",X"83",
		X"81",X"81",X"80",X"80",X"7F",X"7F",X"7D",X"7C",X"7C",X"7C",X"7A",X"7A",X"79",X"79",X"79",X"79",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"76",X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"79",X"79",X"79",X"7A",X"7C",X"7D",X"84",X"90",X"9B",X"A2",
		X"A7",X"A7",X"A5",X"A1",X"9B",X"95",X"8D",X"86",X"7F",X"79",X"71",X"6D",X"67",X"62",X"5F",X"5C",
		X"59",X"58",X"56",X"56",X"56",X"56",X"56",X"58",X"59",X"5B",X"5E",X"5F",X"62",X"65",X"68",X"6B",
		X"6E",X"71",X"74",X"77",X"7A",X"7D",X"80",X"81",X"81",X"80",X"7F",X"7D",X"7D",X"7F",X"80",X"81",
		X"83",X"86",X"89",X"8A",X"8D",X"90",X"93",X"95",X"98",X"99",X"9B",X"9C",X"9E",X"9F",X"9F",X"9F",
		X"9F",X"9F",X"9F",X"9F",X"9E",X"9E",X"9E",X"9C",X"9B",X"99",X"99",X"98",X"9B",X"A2",X"A8",X"AE",
		X"B0",X"B0",X"AD",X"AA",X"A4",X"9E",X"96",X"8F",X"87",X"80",X"79",X"71",X"6B",X"67",X"61",X"5C",
		X"59",X"56",X"53",X"52",X"50",X"50",X"50",X"50",X"50",X"52",X"53",X"56",X"58",X"59",X"5C",X"5F",
		X"61",X"64",X"67",X"6A",X"6D",X"6E",X"71",X"74",X"77",X"79",X"7A",X"7A",X"79",X"76",X"76",X"76",
		X"76",X"77",X"79",X"7C",X"7D",X"80",X"83",X"86",X"89",X"8A",X"8D",X"90",X"92",X"95",X"96",X"98",
		X"99",X"99",X"9B",X"9B",X"9C",X"9B",X"9B",X"9B",X"9B",X"99",X"99",X"98",X"98",X"96",X"95",X"93",
		X"92",X"90",X"8F",X"8D",X"8C",X"8A",X"89",X"87",X"86",X"84",X"84",X"83",X"84",X"89",X"90",X"98",
		X"9E",X"A1",X"A1",X"9F",X"9B",X"96",X"90",X"89",X"81",X"7C",X"74",X"6D",X"67",X"62",X"5C",X"58",
		X"55",X"52",X"4F",X"4D",X"4C",X"4A",X"47",X"43",X"41",X"40",X"40",X"41",X"44",X"49",X"4C",X"52",
		X"56",X"5C",X"62",X"68",X"6D",X"73",X"79",X"7D",X"83",X"87",X"8C",X"90",X"93",X"96",X"99",X"9C",
		X"9E",X"9F",X"A1",X"A2",X"A4",X"A4",X"A4",X"A4",X"A4",X"A4",X"A2",X"A2",X"A1",X"A1",X"A1",X"A5",
		X"AE",X"B4",X"BA",X"BC",X"BA",X"B7",X"B1",X"AB",X"A4",X"9C",X"93",X"8C",X"83",X"7C",X"76",X"6E",
		X"68",X"62",X"5F",X"5B",X"58",X"55",X"53",X"52",X"52",X"52",X"52",X"52",X"53",X"55",X"56",X"58",
		X"59",X"5B",X"5E",X"5C",X"5B",X"5B",X"5B",X"5C",X"5F",X"62",X"65",X"68",X"6D",X"71",X"76",X"7A",
		X"7F",X"83",X"87",X"8C",X"8F",X"92",X"95",X"98",X"9B",X"9C",X"9E",X"9F",X"A1",X"A1",X"A2",X"A2",
		X"A2",X"A2",X"A2",X"A4",X"AA",X"B1",X"B7",X"BC",X"BC",X"BC",X"B9",X"B3",X"AD",X"A7",X"9F",X"98",
		X"8F",X"87",X"80",X"79",X"73",X"6D",X"68",X"64",X"5F",X"5C",X"59",X"56",X"55",X"55",X"53",X"55",
		X"55",X"55",X"56",X"58",X"5B",X"5C",X"5E",X"61",X"62",X"65",X"68",X"6A",X"6B",X"6B",X"6A",X"68",
		X"68",X"6A",X"6A",X"6D",X"6E",X"71",X"76",X"79",X"7C",X"80",X"83",X"86",X"8A",X"8D",X"90",X"92",
		X"95",X"96",X"98",X"9B",X"9B",X"9C",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9C",X"9B",X"99",X"98",
		X"98",X"96",X"95",X"93",X"92",X"90",X"8F",X"8C",X"8A",X"89",X"87",X"86",X"84",X"84",X"86",X"8D",
		X"95",X"9C",X"A2",X"A4",X"A2",X"9F",X"99",X"93",X"8C",X"84",X"7F",X"77",X"70",X"68",X"64",X"5E",
		X"59",X"55",X"52",X"4F",X"4D",X"4C",X"4A",X"4A",X"4C",X"4C",X"4D",X"50",X"52",X"55",X"56",X"58",
		X"56",X"56",X"56",X"56",X"59",X"5C",X"61",X"65",X"6A",X"6E",X"74",X"79",X"7F",X"83",X"87",X"8C",
		X"90",X"95",X"98",X"9B",X"9E",X"A1",X"A4",X"A5",X"A7",X"A8",X"AB",X"B0",X"B9",X"C0",X"C5",X"C8",
		X"C8",X"C5",X"C0",X"BC",X"B6",X"AE",X"A7",X"9E",X"96",X"8F",X"87",X"81",X"7C",X"74",X"70",X"6B",
		X"67",X"62",X"5F",X"5E",X"5B",X"59",X"59",X"59",X"59",X"59",X"5B",X"5B",X"5C",X"5E",X"5F",X"61",
		X"64",X"65",X"67",X"68",X"68",X"67",X"65",X"65",X"65",X"65",X"68",X"6A",X"6D",X"70",X"73",X"77",
		X"7A",X"7F",X"81",X"86",X"89",X"8D",X"8F",X"92",X"95",X"96",X"99",X"9B",X"9C",X"9C",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9C",X"9C",X"9B",X"99",X"99",X"98",X"96",X"93",X"92",X"90",X"8F",X"8D",X"8C",
		X"89",X"87",X"86",X"84",X"83",X"81",X"81",X"81",X"83",X"8A",X"93",X"9B",X"9F",X"A1",X"A1",X"9C",
		X"98",X"92",X"8A",X"84",X"7C",X"76",X"6E",X"68",X"62",X"5C",X"58",X"55",X"52",X"4F",X"4D",X"4D",
		X"4C",X"4C",X"4D",X"4D",X"4F",X"50",X"53",X"55",X"58",X"5B",X"5F",X"62",X"65",X"6A",X"6D",X"70",
		X"74",X"77",X"7A",X"7D",X"80",X"83",X"84",X"87",X"89",X"8A",X"8D",X"8F",X"8F",X"90",X"92",X"92",
		X"93",X"93",X"92",X"8D",X"89",X"86",X"84",X"83",X"81",X"83",X"83",X"83",X"84",X"86",X"87",X"89",
		X"8A",X"8C",X"8D",X"8F",X"90",X"90",X"92",X"92",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"93",
		X"92",X"90",X"90",X"8F",X"8D",X"8D",X"8C",X"8A",X"89",X"89",X"87",X"86",X"84",X"83",X"83",X"81",
		X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"81",X"89",X"92",X"99",X"9E",X"A1",X"9F",X"9C",X"98",X"93",
		X"8C",X"86",X"7F",X"77",X"71",X"6B",X"65",X"61",X"5C",X"58",X"55",X"53",X"50",X"4F",X"4F",X"4F",
		X"4F",X"50",X"52",X"53",X"55",X"58",X"59",X"5C",X"5F",X"62",X"65",X"68",X"6B",X"6E",X"70",X"73",
		X"73",X"71",X"70",X"70",X"71",X"73",X"74",X"77",X"7A",X"7F",X"81",X"84",X"89",X"8C",X"8F",X"93",
		X"96",X"98",X"9B",X"9C",X"9E",X"A1",X"A1",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A2",X"A1",
		X"A1",X"A5",X"AB",X"B3",X"B9",X"BA",X"BA",X"B7",X"B3",X"AD",X"A5",X"9F",X"96",X"8F",X"87",X"80",
		X"79",X"71",X"6B",X"65",X"61",X"5E",X"59",X"56",X"55",X"53",X"52",X"50",X"50",X"50",X"52",X"50",
		X"4F",X"4C",X"4A",X"4A",X"4C",X"4F",X"52",X"55",X"59",X"5E",X"62",X"68",X"6D",X"71",X"77",X"7C",
		X"80",X"84",X"87",X"8C",X"8F",X"92",X"95",X"98",X"99",X"9B",X"9C",X"9E",X"9E",X"9F",X"9F",X"9F",
		X"9F",X"9F",X"9E",X"9E",X"9E",X"9C",X"9F",X"A7",X"AE",X"B4",X"B6",X"B7",X"B6",X"B1",X"AB",X"A5",
		X"9E",X"96",X"8D",X"86",X"7F",X"77",X"70",X"6A",X"65",X"5F",X"5B",X"58",X"55",X"53",X"52",X"50",
		X"50",X"50",X"52",X"52",X"53",X"55",X"56",X"59",X"5C",X"5E",X"61",X"64",X"67",X"6A",X"6D",X"70",
		X"73",X"76",X"77",X"7A",X"7C",X"7D",X"7C",X"7A",X"79",X"79",X"79",X"7A",X"7C",X"7D",X"7F",X"81",
		X"84",X"87",X"89",X"8C",X"8F",X"90",X"93",X"95",X"98",X"99",X"99",X"9B",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9C",X"9B",X"9B",X"99",X"99",X"98",X"98",X"96",X"98",X"9E",X"A5",X"AB",X"AE",X"B0",X"AE",
		X"AB",X"A7",X"A1",X"99",X"92",X"8A",X"81",X"7C",X"74",X"6D",X"67",X"62",X"5E",X"59",X"56",X"53",
		X"52",X"50",X"4F",X"4F",X"4F",X"4F",X"50",X"52",X"53",X"56",X"58",X"5B",X"5E",X"61",X"64",X"67",
		X"6A",X"6D",X"70",X"73",X"76",X"77",X"7A",X"7D",X"7F",X"81",X"83",X"84",X"87",X"87",X"89",X"8A",
		X"8C",X"8A",X"87",X"84",X"81",X"80",X"80",X"80",X"80",X"81",X"83",X"84",X"86",X"87",X"89",X"8A",
		X"8D",X"8F",X"90",X"92",X"93",X"93",X"95",X"95",X"96",X"96",X"96",X"96",X"95",X"95",X"95",X"93",
		X"93",X"92",X"92",X"92",X"90",X"8F",X"8F",X"8F",X"92",X"99",X"A1",X"A5",X"A7",X"A7",X"A5",X"A1",
		X"9C",X"96",X"8F",X"87",X"81",X"7A",X"74",X"6D",X"67",X"62",X"5E",X"5B",X"56",X"53",X"52",X"50",
		X"50",X"50",X"50",X"52",X"52",X"53",X"55",X"58",X"59",X"5C",X"5F",X"62",X"64",X"67",X"6A",X"6D",
		X"70",X"73",X"76",X"79",X"7A",X"7D",X"80",X"81",X"83",X"84",X"86",X"87",X"89",X"8A",X"8C",X"8A",
		X"87",X"84",X"81",X"80",X"7F",X"7F",X"7F",X"80",X"81",X"83",X"84",X"86",X"87",X"8A",X"8C",X"8D",
		X"8F",X"90",X"92",X"93",X"95",X"95",X"96",X"96",X"96",X"96",X"96",X"96",X"96",X"96",X"96",X"95",
		X"95",X"95",X"95",X"96",X"9E",X"A4",X"AA",X"AD",X"AD",X"AB",X"A8",X"A2",X"9C",X"96",X"8F",X"87",
		X"80",X"7A",X"73",X"6D",X"67",X"62",X"5E",X"5B",X"58",X"55",X"53",X"52",X"52",X"52",X"52",X"52",
		X"53",X"55",X"56",X"59",X"5B",X"5E",X"5F",X"62",X"65",X"68",X"6A",X"6D",X"70",X"73",X"74",X"77",
		X"79",X"7A",X"7A",X"79",X"77",X"76",X"74",X"76",X"77",X"79",X"7A",X"7C",X"7F",X"81",X"84",X"87",
		X"8A",X"8D",X"90",X"92",X"95",X"96",X"98",X"99",X"9B",X"9C",X"9C",X"9E",X"9E",X"9E",X"9E",X"9C",
		X"9C",X"9C",X"9B",X"9B",X"99",X"98",X"96",X"95",X"93",X"92",X"90",X"8F",X"8D",X"8C",X"8A",X"89",
		X"86",X"86",X"84",X"84",X"89",X"8F",X"95",X"99",X"9B",X"99",X"96",X"93",X"8D",X"87",X"81",X"7C",
		X"76",X"70",X"6A",X"65",X"5F",X"5C",X"59",X"56",X"53",X"52",X"50",X"50",X"50",X"50",X"52",X"53",
		X"55",X"58",X"59",X"5C",X"5F",X"61",X"64",X"67",X"6A",X"6B",X"6D",X"6B",X"6B",X"6A",X"6B",X"6B",
		X"6E",X"70",X"73",X"77",X"7A",X"7D",X"81",X"84",X"89",X"8C",X"90",X"93",X"96",X"99",X"9B",X"9E",
		X"9F",X"A1",X"A1",X"A2",X"A2",X"A4",X"A4",X"A4",X"A4",X"A4",X"A2",X"A1",X"9F",X"9E",X"9C",X"9B",
		X"99",X"98",X"96",X"95",X"93",X"92",X"92",X"96",X"9C",X"A1",X"A2",X"A2",X"A1",X"9E",X"98",X"92",
		X"8C",X"86",X"7F",X"79",X"71",X"6B",X"67",X"61",X"5E",X"59",X"56",X"53",X"52",X"50",X"4F",X"4D",
		X"4A",X"46",X"43",X"43",X"43",X"46",X"49",X"4C",X"50",X"55",X"59",X"5F",X"65",X"6A",X"70",X"76",
		X"7A",X"80",X"84",X"89",X"8D",X"90",X"95",X"98",X"9B",X"9C",X"9E",X"9F",X"A1",X"A2",X"A2",X"A4",
		X"A4",X"A4",X"A4",X"A7",X"AE",X"B4",X"B7",X"B9",X"B7",X"B4",X"B0",X"AB",X"A4",X"9E",X"96",X"8F",
		X"87",X"80",X"79",X"73",X"6D",X"68",X"64",X"61",X"5E",X"5B",X"59",X"58",X"58",X"56",X"56",X"58",
		X"59",X"59",X"5B",X"5E",X"5F",X"62",X"64",X"67",X"68",X"6B",X"6E",X"70",X"73",X"76",X"79",X"7A",
		X"7D",X"7F",X"80",X"83",X"84",X"84",X"86",X"86",X"83",X"80",X"7D",X"7D",X"7C",X"7C",X"7D",X"7D",
		X"7F",X"80",X"83",X"84",X"86",X"89",X"8A",X"8D",X"8F",X"90",X"92",X"93",X"95",X"96",X"96",X"96",
		X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"98",X"99",X"9E",X"A5",X"AA",X"AD",X"AD",X"AA",X"A7",
		X"A2",X"9C",X"96",X"8F",X"89",X"81",X"7C",X"76",X"70",X"6A",X"65",X"61",X"5E",X"5B",X"58",X"56",
		X"56",X"55",X"55",X"55",X"55",X"56",X"58",X"59",X"5B",X"5E",X"5F",X"62",X"64",X"67",X"6A",X"6B",
		X"6E",X"71",X"73",X"76",X"77",X"7A",X"7C",X"7C",X"79",X"77",X"76",X"76",X"76",X"77",X"79",X"7A",
		X"7D",X"7F",X"81",X"84",X"87",X"8A",X"8C",X"8F",X"92",X"93",X"96",X"98",X"99",X"9B",X"9C",X"9C",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9C",X"9C",X"9B",X"9B",X"99",X"99",X"9E",X"A4",X"A8",X"AA",X"AA",
		X"A8",X"A5",X"A1",X"9B",X"93",X"8D",X"87",X"80",X"7A",X"74",X"6E",X"68",X"64",X"5F",X"5C",X"59",
		X"58",X"56",X"55",X"55",X"55",X"55",X"56",X"56",X"58",X"59",X"5B",X"5C",X"5F",X"61",X"64",X"67",
		X"6A",X"6B",X"6E",X"71",X"73",X"76",X"79",X"7A",X"7C",X"7D",X"7C",X"79",X"77",X"77",X"77",X"77",
		X"79",X"7A",X"7C",X"7F",X"80",X"83",X"86",X"89",X"8C",X"8F",X"90",X"93",X"95",X"98",X"98",X"9B",
		X"9C",X"9C",X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"9C",X"9C",X"9B",X"99",X"98",X"96",X"95",X"93",
		X"90",X"8F",X"8D",X"8C",X"8A",X"8A",X"8F",X"95",X"98",X"99",X"99",X"98",X"93",X"90",X"8A",X"84",
		X"80",X"7A",X"74",X"70",X"6A",X"65",X"61",X"5E",X"5C",X"59",X"58",X"56",X"56",X"55",X"55",X"55",
		X"56",X"55",X"52",X"50",X"4F",X"4F",X"50",X"53",X"56",X"5B",X"5F",X"64",X"68",X"6E",X"73",X"79",
		X"7D",X"81",X"86",X"8C",X"8F",X"93",X"96",X"99",X"9C",X"9F",X"A1",X"A2",X"A4",X"A5",X"A7",X"AA",
		X"B0",X"B4",X"B9",X"BA",X"BA",X"B7",X"B4",X"AE",X"A8",X"A2",X"9C",X"95",X"8D",X"87",X"81",X"7C",
		X"76",X"71",X"6D",X"68",X"65",X"62",X"61",X"5F",X"5E",X"5C",X"5C",X"5C",X"5C",X"5E",X"5F",X"61",
		X"61",X"62",X"64",X"67",X"68",X"6A",X"6D",X"6E",X"70",X"71",X"73",X"74",X"71",X"70",X"6E",X"6E",
		X"6E",X"70",X"71",X"74",X"77",X"7A",X"7D",X"81",X"84",X"87",X"8C",X"8F",X"90",X"93",X"96",X"98",
		X"9B",X"9C",X"9E",X"9F",X"9F",X"A1",X"A2",X"A8",X"AE",X"B3",X"B4",X"B6",X"B4",X"B0",X"AB",X"A7",
		X"A1",X"9B",X"93",X"8D",X"87",X"81",X"7A",X"76",X"71",X"6D",X"68",X"65",X"62",X"5F",X"5E",X"5C",
		X"5C",X"5B",X"5B",X"5B",X"5C",X"5C",X"5E",X"5F",X"61",X"62",X"64",X"67",X"68",X"6A",X"6D",X"6E",
		X"71",X"73",X"74",X"76",X"77",X"77",X"74",X"73",X"71",X"71",X"71",X"73",X"74",X"76",X"79",X"7C",
		X"7F",X"81",X"84",X"87",X"8A",X"8D",X"90",X"93",X"95",X"98",X"99",X"9C",X"9C",X"9E",X"9E",X"9E",
		X"9E",X"9E",X"9E",X"9C",X"9B",X"99",X"98",X"96",X"95",X"93",X"92",X"8F",X"8D",X"8C",X"8A",X"87",
		X"86",X"83",X"81",X"80",X"7F",X"7D",X"7C",X"79",X"79",X"77",X"76",X"76",X"76",X"76",X"77",X"7C",
		X"81",X"86",X"89",X"89",X"89",X"87",X"84",X"81",X"7F",X"7A",X"77",X"73",X"70",X"6D",X"6A",X"67",
		X"64",X"62",X"61",X"61",X"61",X"5F",X"61",X"61",X"61",X"62",X"64",X"65",X"67",X"6A",X"6B",X"6D",
		X"70",X"73",X"74",X"76",X"79",X"7A",X"7C",X"7F",X"80",X"81",X"83",X"84",X"86",X"87",X"89",X"89",
		X"8A",X"8A",X"8C",X"8C",X"8C",X"8D",X"8D",X"8F",X"8F",X"8F",X"8D",X"8D",X"8D",X"8D",X"8C",X"8C",
		X"8A",X"86",X"81",X"7D",X"7A",X"79",X"77",X"77",X"77",X"77",X"79",X"7A",X"7C",X"7F",X"81",X"83",
		X"86",X"87",X"8A",X"8C",X"8D",X"90",X"92",X"92",X"93",X"93",X"93",X"93",X"93",X"93",X"93",X"92",
		X"90",X"90",X"8F",X"8D",X"8C",X"8A",X"89",X"87",X"86",X"84",X"83",X"81",X"80",X"7F",X"7D",X"7C",
		X"7A",X"79",X"79",X"77",X"77",X"76",X"76",X"77",X"7C",X"80",X"84",X"87",X"89",X"89",X"87",X"84",
		X"81",X"7F",X"7A",X"77",X"73",X"70",X"6D",X"6A",X"67",X"65",X"64",X"62",X"61",X"61",X"61",X"61",
		X"61",X"61",X"62",X"64",X"65",X"67",X"68",X"6A",X"6D",X"70",X"71",X"73",X"76",X"79",X"7A",X"7C",
		X"7F",X"80",X"81",X"83",X"84",X"86",X"87",X"89",X"89",X"89",X"86",X"81",X"80",X"7F",X"7D",X"7D",
		X"7D",X"7F",X"80",X"81",X"84",X"86",X"89",X"8C",X"8D",X"90",X"92",X"95",X"96",X"98",X"99",X"99",
		X"9B",X"9B",X"9B",X"9B",X"99",X"99",X"98",X"96",X"95",X"93",X"93",X"90",X"8F",X"8D",X"8A",X"89",
		X"87",X"86",X"84",X"83",X"81",X"80",X"7F",X"7D",X"7F",X"83",X"86",X"89",X"8A",X"8A",X"89",X"86",
		X"83",X"80",X"7C",X"79",X"74",X"71",X"6E",X"6A",X"67",X"65",X"62",X"61",X"5F",X"5F",X"5F",X"5F",
		X"5F",X"5F",X"61",X"61",X"62",X"64",X"67",X"68",X"6A",X"6B",X"6D",X"70",X"71",X"73",X"74",X"74",
		X"71",X"71",X"70",X"70",X"70",X"73",X"74",X"77",X"7A",X"7D",X"81",X"84",X"87",X"8C",X"8F",X"92",
		X"95",X"98",X"99",X"9B",X"9E",X"9E",X"9F",X"9F",X"9F",X"9F",X"9F",X"9E",X"9E",X"9C",X"9B",X"99",
		X"98",X"96",X"93",X"92",X"90",X"8D",X"8C",X"89",X"87",X"86",X"84",X"83",X"80",X"80",X"7D",X"7C",
		X"7C",X"7A",X"79",X"77",X"77",X"76",X"76",X"74",X"74",X"74",X"74",X"74",X"74",X"74",X"77",X"7C",
		X"81",X"84",X"87",X"89",X"87",X"87",X"84",X"83",X"80",X"7D",X"7A",X"76",X"73",X"71",X"6E",X"6D",
		X"6B",X"6A",X"68",X"68",X"67",X"67",X"67",X"67",X"68",X"68",X"65",X"62",X"5F",X"5E",X"5F",X"5F",
		X"62",X"64",X"68",X"6B",X"70",X"74",X"79",X"7D",X"81",X"86",X"8A",X"8D",X"90",X"95",X"96",X"99",
		X"9B",X"9C",X"9E",X"9F",X"9F",X"9F",X"9F",X"A1",X"A2",X"A5",X"AA",X"AB",X"AB",X"AB",X"A8",X"A5",
		X"A1",X"9C",X"96",X"92",X"8C",X"87",X"81",X"7D",X"79",X"76",X"73",X"70",X"6D",X"6A",X"68",X"67",
		X"65",X"65",X"65",X"64",X"65",X"65",X"65",X"67",X"67",X"68",X"6A",X"6B",X"6D",X"6E",X"70",X"71",
		X"73",X"74",X"76",X"77",X"76",X"74",X"71",X"70",X"70",X"70",X"71",X"73",X"74",X"77",X"7A",X"7D",
		X"80",X"83",X"86",X"89",X"8C",X"8F",X"92",X"93",X"95",X"96",X"98",X"99",X"99",X"99",X"99",X"98",
		X"98",X"96",X"96",X"95",X"93",X"92",X"90",X"8F",X"8D",X"8C",X"8A",X"89",X"86",X"84",X"84",X"83",
		X"81",X"84",X"87",X"8A",X"8C",X"8C",X"8C",X"8A",X"87",X"84",X"80",X"7D",X"79",X"76",X"73",X"70",
		X"6D",X"6A",X"68",X"67",X"65",X"64",X"64",X"64",X"64",X"64",X"64",X"65",X"65",X"67",X"68",X"6A",
		X"6B",X"6D",X"6E",X"70",X"71",X"70",X"6D",X"6B",X"6A",X"6B",X"6D",X"6E",X"71",X"74",X"77",X"7C",
		X"7F",X"81",X"86",X"89",X"8C",X"8F",X"92",X"95",X"96",X"98",X"99",X"9B",X"9C",X"9C",X"9C",X"9C",
		X"9C",X"9B",X"99",X"99",X"98",X"96",X"96",X"95",X"93",X"95",X"98",X"99",X"99",X"99",X"98",X"96",
		X"93",X"8F",X"8C",X"87",X"83",X"7F",X"7A",X"77",X"73",X"70",X"6D",X"6A",X"68",X"65",X"65",X"64",
		X"64",X"62",X"62",X"62",X"64",X"64",X"65",X"67",X"67",X"68",X"6A",X"6D",X"6E",X"70",X"71",X"73",
		X"74",X"76",X"76",X"74",X"73",X"71",X"70",X"70",X"71",X"73",X"76",X"79",X"7C",X"7F",X"81",X"84",
		X"87",X"8C",X"8D",X"90",X"93",X"95",X"96",X"98",X"99",X"99",X"99",X"99",X"99",X"99",X"98",X"98",
		X"96",X"95",X"93",X"92",X"90",X"8F",X"8D",X"8C",X"89",X"87",X"86",X"84",X"83",X"81",X"80",X"7F",
		X"7F",X"7D",X"7C",X"7A",X"7A",X"79",X"79",X"77",X"77",X"77",X"76",X"76",X"76",X"76",X"76",X"76",
		X"76",X"76",X"76",X"76",X"77",X"7A",X"7F",X"83",X"86",X"87",X"89",X"89",X"87",X"86",X"84",X"81",
		X"80",X"7D",X"7C",X"79",X"77",X"74",X"73",X"71",X"70",X"70",X"6E",X"6E",X"6E",X"6E",X"6E",X"70",
		X"70",X"70",X"71",X"73",X"73",X"74",X"74",X"76",X"77",X"79",X"7A",X"7C",X"7D",X"7D",X"7F",X"80",
		X"80",X"81",X"83",X"83",X"83",X"84",X"84",X"86",X"86",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"89",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"86",X"86",X"84",X"80",X"7C",X"79",X"77",X"76",
		X"76",X"76",X"77",X"79",X"7A",X"7D",X"7F",X"80",X"83",X"86",X"87",X"89",X"8A",X"8C",X"8D",X"8F",
		X"8F",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8F",X"8D",X"8C",X"8C",X"8A",X"89",X"87",X"86",X"86",
		X"83",X"83",X"81",X"80",X"7F",X"7D",X"7D",X"7C",X"7A",X"7A",X"79",X"79",X"77",X"76",X"76",X"76",
		X"76",X"76",X"74",X"74",X"76",X"76",X"76",X"79",X"7C",X"80",X"83",X"84",X"84",X"84",X"84",X"83",
		X"80",X"7F",X"7D",X"7A",X"79",X"77",X"74",X"73",X"71",X"70",X"70",X"6E",X"6E",X"6E",X"6E",X"6E",
		X"6E",X"6E",X"70",X"70",X"71",X"73",X"74",X"76",X"77",X"77",X"79",X"7A",X"7C",X"7D",X"7D",X"7F",
		X"7F",X"7D",X"7A",X"79",X"77",X"77",X"79",X"7A",X"7C",X"7F",X"80",X"83",X"86",X"89",X"8C",X"8D",
		X"8F",X"92",X"93",X"95",X"95",X"96",X"96",X"96",X"96",X"96",X"96",X"95",X"95",X"93",X"92",X"92",
		X"90",X"8F",X"8C",X"8A",X"89",X"87",X"86",X"86",X"84",X"83",X"81",X"80",X"80",X"81",X"84",X"86",
		X"87",X"87",X"87",X"86",X"83",X"81",X"7F",X"7C",X"79",X"76",X"73",X"71",X"6E",X"6D",X"6B",X"6A",
		X"6A",X"68",X"68",X"68",X"67",X"68",X"68",X"68",X"6A",X"6B",X"6D",X"6E",X"70",X"71",X"73",X"74",
		X"76",X"77",X"77",X"7A",X"7A",X"7C",X"7D",X"7F",X"7F",X"7D",X"7A",X"79",X"79",X"79",X"79",X"7A",
		X"7C",X"7F",X"80",X"83",X"86",X"87",X"8A",X"8C",X"8F",X"90",X"92",X"92",X"93",X"95",X"95",X"95",
		X"95",X"95",X"95",X"93",X"93",X"92",X"90",X"90",X"8F",X"8D",X"8C",X"8A",X"89",X"87",X"86",X"86",
		X"84",X"83",X"81",X"81",X"81",X"83",X"86",X"87",X"89",X"89",X"87",X"86",X"83",X"81",X"7F",X"7C",
		X"79",X"77",X"74",X"73",X"70",X"6E",X"6D",X"6B",X"6B",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",X"6A",
		X"6B",X"6D",X"6D",X"6E",X"70",X"70",X"71",X"73",X"74",X"76",X"77",X"79",X"79",X"7A",X"79",X"76",
		X"74",X"74",X"74",X"76",X"77",X"7A",X"7D",X"7F",X"81",X"84",X"87",X"89",X"8C",X"8F",X"90",X"92",
		X"93",X"93",X"95",X"95",X"95",X"95",X"95",X"95",X"95",X"93",X"92",X"92",X"90",X"8F",X"8D",X"8C",
		X"8A",X"89",X"89",X"87",X"86",X"84",X"83",X"81",X"80",X"80",X"7F",X"7F",X"7D",X"7C",X"7C",X"7D",
		X"7F",X"81",X"83",X"83",X"83",X"83",X"81",X"80",X"7F",X"7C",X"7A",X"79",X"76",X"74",X"73",X"71",
		X"70",X"70",X"70",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"70",X"70",X"70",X"70",X"6E",X"6D",
		X"6B",X"6B",X"6D",X"6E",X"70",X"73",X"76",X"77",X"7A",X"7D",X"80",X"83",X"86",X"87",X"8A",X"8C",
		X"8D",X"8F",X"90",X"92",X"92",X"92",X"93",X"92",X"92",X"92",X"92",X"90",X"90",X"8F",X"8F",X"8D",
		X"8C",X"8A",X"8A",X"89",X"87",X"86",X"84",X"84",X"83",X"81",X"81",X"80",X"80",X"7F",X"7F",X"80",
		X"80",X"81",X"83",X"83",X"83",X"81",X"80",X"80",X"7F",X"7D",X"7C",X"7A",X"79",X"77",X"76",X"74",
		X"73",X"73",X"73",X"71",X"71",X"71",X"71",X"71",X"71",X"73",X"73",X"74",X"74",X"76",X"76",X"76",
		X"76",X"74",X"73",X"73",X"73",X"73",X"74",X"76",X"77",X"79",X"7A",X"7D",X"7F",X"81",X"83",X"84",
		X"87",X"89",X"8A",X"8C",X"8D",X"8D",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8D",X"8D",X"8D",
		X"8C",X"8C",X"8A",X"89",X"87",X"87",X"86",X"86",X"84",X"83",X"81",X"81",X"80",X"80",X"7F",X"7F",
		X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7D",
		X"80",X"83",X"84",X"86",X"86",X"86",X"84",X"84",X"83",X"80",X"7F",X"7D",X"7C",X"7A",X"79",X"77",
		X"76",X"76",X"74",X"74",X"74",X"74",X"73",X"73",X"73",X"73",X"74",X"74",X"74",X"76",X"76",X"77",
		X"77",X"79",X"79",X"7A",X"7C",X"7C",X"7D",X"7D",X"7D",X"7C",X"7A",X"79",X"77",X"77",X"79",X"7A",
		X"7A",X"7D",X"7F",X"81",X"83",X"84",X"87",X"89",X"8A",X"8C",X"8D",X"8F",X"8F",X"8F",X"90",X"90",
		X"90",X"90",X"8F",X"8F",X"8F",X"8D",X"8D",X"8C",X"8C",X"8A",X"89",X"89",X"87",X"86",X"86",X"84",
		X"84",X"83",X"84",X"86",X"87",X"87",X"87",X"87",X"86",X"84",X"83",X"81",X"7F",X"7D",X"7A",X"79",
		X"76",X"74",X"73",X"71",X"71",X"70",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"70",
		X"6E",X"6D",X"6B",X"6B",X"6B",X"6B",X"6D",X"70",X"71",X"74",X"77",X"79",X"7C",X"7F",X"81",X"83",
		X"86",X"87",X"89",X"8A",X"8C",X"8D",X"8F",X"8F",X"90",X"90",X"90",X"90",X"90",X"8F",X"8F",X"8D",
		X"8D",X"8D",X"8C",X"8C",X"8A",X"89",X"89",X"8A",X"8C",X"8D",X"8D",X"8D",X"8C",X"8A",X"89",X"87",
		X"84",X"83",X"80",X"7D",X"7C",X"79",X"77",X"76",X"74",X"73",X"71",X"71",X"70",X"70",X"70",X"70",
		X"70",X"70",X"70",X"70",X"71",X"71",X"73",X"74",X"74",X"76",X"76",X"77",X"79",X"79",X"7A",X"7A",
		X"7A",X"79",X"77",X"76",X"76",X"76",X"77",X"79",X"7A",X"7D",X"7F",X"80",X"83",X"84",X"86",X"89",
		X"8A",X"8A",X"8C",X"8D",X"8D",X"8D",X"8F",X"8F",X"8F",X"8F",X"8F",X"8F",X"8D",X"8D",X"8D",X"8C",
		X"8C",X"8A",X"89",X"89",X"89",X"8A",X"8C",X"8C",X"8C",X"8C",X"8A",X"89",X"86",X"84",X"83",X"80",
		X"7D",X"7C",X"79",X"77",X"76",X"74",X"73",X"71",X"71",X"70",X"70",X"6E",X"6E",X"6E",X"6E",X"70",
		X"70",X"71",X"71",X"73",X"73",X"74",X"74",X"76",X"77",X"79",X"79",X"7A",X"7A",X"7C",X"7C",X"7D",
		X"7F",X"7F",X"7F",X"7F",X"7D",X"7C",X"7A",X"7A",X"7A",X"7A",X"7C",X"7D",X"7F",X"80",X"81",X"83",
		X"84",X"86",X"87",X"89",X"8A",X"8A",X"8A",X"8C",X"8C",X"8D",X"8D",X"8D",X"8C",X"8C",X"8C",X"8A",
		X"8A",X"8A",X"89",X"89",X"87",X"86",X"86",X"84",X"83",X"83",X"81",X"81",X"80",X"80",X"7F",X"7F",
		X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7F",X"80",X"81",X"83",X"81",X"81",X"81",
		X"80",X"7F",X"7D",X"7D",X"7C",X"7A",X"79",X"77",X"76",X"76",X"74",X"74",X"74",X"74",X"74",X"74",
		X"74",X"74",X"74",X"76",X"76",X"76",X"77",X"77",X"79",X"79",X"7A",X"7A",X"7C",X"7C",X"7D",X"7D",
		X"7F",X"7F",X"80",X"80",X"7F",X"7D",X"7C",X"7A",X"7A",X"7A",X"7C",X"7C",X"7D",X"7F",X"80",X"81",
		X"83",X"84",X"86",X"87",X"89",X"89",X"8A",X"8A",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",X"8C",
		X"8A",X"8A",X"89",X"89",X"87",X"87",X"86",X"86",X"84",X"84",X"83",X"83",X"81",X"81",X"80",X"80",
		X"7F",X"7F",X"7F",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7C",X"7D",X"7F",X"81",X"81",X"83",X"83",X"81",X"81",X"80",X"80",X"7F",X"7D",X"7D",X"7C",X"7A",
		X"7A",X"79",X"77",X"77",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"76",X"77",X"77",X"77",
		X"79",X"79",X"79",X"7A",X"7A",X"7C",X"7C",X"7D",X"7D",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",
		X"83",X"83",X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"83",X"83",X"83",X"83",X"80",X"7F",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7F",X"7F",X"80",
		X"81",X"83",X"83",X"84",X"86",X"86",X"86",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"86",
		X"86",X"84",X"84",X"84",X"83",X"83",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7D",X"7D",
		X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",
		X"7C",X"7D",X"80",X"81",X"81",X"83",X"83",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7D",X"7C",X"7C",
		X"7A",X"79",X"79",X"79",X"77",X"77",X"77",X"77",X"77",X"77",X"79",X"79",X"79",X"79",X"7A",X"7A",
		X"7A",X"7A",X"7A",X"79",X"77",X"77",X"77",X"79",X"79",X"7A",X"7C",X"7D",X"7F",X"80",X"81",X"83",
		X"84",X"86",X"87",X"89",X"89",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"8A",X"89",
		X"89",X"89",X"89",X"87",X"86",X"86",X"86",X"84",X"84",X"86",X"86",X"87",X"87",X"87",X"86",X"84",
		X"83",X"83",X"80",X"7F",X"7D",X"7C",X"7A",X"79",X"79",X"77",X"76",X"76",X"74",X"74",X"74",X"74",
		X"74",X"74",X"74",X"74",X"74",X"74",X"76",X"77",X"77",X"79",X"79",X"79",X"7A",X"7A",X"7C",X"7C",
		X"7C",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7F",
		X"7F",X"80",X"81",X"81",X"83",X"84",X"86",X"86",X"87",X"87",X"89",X"89",X"89",X"89",X"89",X"89",
		X"89",X"89",X"89",X"89",X"8A",X"8C",X"8C",X"8C",X"8A",X"8A",X"89",X"87",X"86",X"84",X"83",X"81",
		X"80",X"7F",X"7D",X"7C",X"7A",X"79",X"79",X"77",X"77",X"76",X"76",X"76",X"76",X"76",X"76",X"76",
		X"76",X"76",X"76",X"77",X"77",X"77",X"77",X"79",X"79",X"7A",X"7A",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7A",X"7A",X"79",X"79",X"79",X"7A",X"7C",X"7C",X"7D",X"7F",X"80",X"81",X"83",X"83",X"84",X"84",
		X"86",X"86",X"87",X"87",X"87",X"89",X"89",X"89",X"89",X"87",X"87",X"87",X"87",X"86",X"86",X"86",
		X"86",X"84",X"84",X"83",X"83",X"83",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7D",X"7F",X"80",X"80",X"81",X"81",X"83",X"81",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7D",
		X"7D",X"7C",X"7C",X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",
		X"7A",X"7A",X"79",X"79",X"77",X"79",X"79",X"79",X"7A",X"7C",X"7C",X"7D",X"7F",X"80",X"81",X"83",
		X"83",X"84",X"84",X"86",X"86",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"89",X"89",X"8A",X"89",X"89",X"89",X"87",X"86",X"84",X"83",X"81",X"80",X"80",X"7F",X"7D",X"7C",
		X"7C",X"7A",X"7A",X"79",X"79",X"79",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"79",X"79",X"79",
		X"79",X"79",X"7A",X"79",X"79",X"77",X"77",X"77",X"79",X"79",X"7A",X"7A",X"7C",X"7D",X"7F",X"80",
		X"80",X"81",X"83",X"83",X"84",X"84",X"86",X"86",X"86",X"86",X"87",X"87",X"87",X"86",X"86",X"86",
		X"86",X"86",X"86",X"84",X"84",X"84",X"83",X"83",X"83",X"81",X"81",X"81",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"7F",X"7F",
		X"7D",X"7D",X"7C",X"7C",X"7A",X"7A",X"7A",X"7A",X"79",X"79",X"79",X"79",X"79",X"79",X"79",X"79",
		X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7D",X"7D",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7F",X"7F",X"80",X"80",X"81",X"83",X"83",X"84",X"84",X"84",
		X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"86",X"84",X"84",X"84",X"83",
		X"83",X"83",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7D",X"7D",X"7C",X"7C",X"7C",X"7A",X"7A",X"7A",X"7A",X"7C",X"7A",X"7A",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"80",
		X"80",X"80",X"81",X"81",X"83",X"83",X"83",X"83",X"83",X"84",X"84",X"84",X"84",X"84",X"84",X"84",
		X"84",X"84",X"84",X"83",X"83",X"83",X"83",X"83",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"80",X"80",X"80",X"81",X"81",X"83",X"83",X"83",X"83",X"84",
		X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"84",X"83",X"83",X"83",X"83",X"83",X"83",X"84",
		X"84",X"83",X"83",X"83",X"81",X"81",X"81",X"80",X"80",X"7F",X"7F",X"7D",X"7D",X"7D",X"7C",X"7C",
		X"7C",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7A",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7A",X"7A",X"7C",X"7C",X"7C",X"7D",X"7D",X"7F",X"7F",X"7F",X"80",X"80",
		X"81",X"81",X"81",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",
		X"83",X"83",X"83",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7F",X"7F",X"7F",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",
		X"80",X"81",X"81",X"81",X"81",X"83",X"81",X"83",X"83",X"83",X"83",X"81",X"83",X"83",X"83",X"83",
		X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"81",X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",
		X"7F",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"81",
		X"81",X"81",X"81",X"81",X"81",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"83",X"81",X"81",
		X"81",X"81",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7C",X"7C",X"7C",X"7C",X"7D",X"7D",
		X"7D",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"80",X"81",X"81",X"81",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7D",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",
		X"80",X"80",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",X"81",
		X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7D",X"7D",X"7D",
		X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"81",X"81",X"81",X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7D",X"7F",X"7D",X"7D",X"7D",
		X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"81",X"81",X"81",
		X"81",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7D",X"7F",X"7D",X"7F",X"7D",X"7D",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",
		X"7F",X"7F",X"80",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"7F",X"80",X"7F",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",
		X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",
		X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",
		X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"82",
		X"7C",X"7C",X"80",X"87",X"87",X"7C",X"80",X"8B",X"82",X"7C",X"82",X"87",X"82",X"77",X"69",X"7C",
		X"90",X"B1",X"DB",X"D7",X"B6",X"95",X"6E",X"7C",X"95",X"BA",X"DB",X"BF",X"9E",X"82",X"A3",X"B1",
		X"9E",X"B6",X"B6",X"A7",X"87",X"87",X"A7",X"C8",X"BF",X"90",X"7C",X"82",X"82",X"82",X"80",X"7C",
		X"82",X"82",X"80",X"7C",X"82",X"87",X"99",X"99",X"82",X"69",X"43",X"56",X"7C",X"99",X"B6",X"95",
		X"77",X"51",X"43",X"69",X"82",X"A7",X"AC",X"82",X"69",X"43",X"51",X"77",X"90",X"B1",X"99",X"77",
		X"56",X"3F",X"64",X"80",X"A3",X"AC",X"87",X"69",X"48",X"27",X"31",X"51",X"72",X"90",X"80",X"60",
		X"43",X"60",X"82",X"A3",X"B6",X"8B",X"72",X"4D",X"48",X"72",X"8B",X"B1",X"9E",X"80",X"60",X"43",
		X"5B",X"80",X"95",X"72",X"64",X"87",X"90",X"69",X"6E",X"8B",X"AC",X"D2",X"BF",X"9E",X"80",X"90",
		X"B1",X"D2",X"E5",X"C4",X"A7",X"80",X"7C",X"95",X"BA",X"BA",X"90",X"72",X"51",X"35",X"43",X"64",
		X"82",X"69",X"51",X"69",X"51",X"4D",X"5B",X"7C",X"82",X"5B",X"60",X"64",X"4D",X"31",X"3F",X"64",
		X"7C",X"6E",X"48",X"31",X"51",X"77",X"90",X"B6",X"BA",X"99",X"7C",X"56",X"5B",X"80",X"9E",X"90",
		X"69",X"4D",X"2C",X"14",X"31",X"51",X"77",X"82",X"69",X"43",X"3F",X"69",X"82",X"A7",X"9E",X"77",
		X"5B",X"69",X"60",X"4D",X"60",X"6E",X"5B",X"51",X"64",X"7C",X"A7",X"A3",X"87",X"64",X"69",X"8B",
		X"80",X"82",X"99",X"87",X"7C",X"4D",X"3F",X"5B",X"80",X"87",X"80",X"87",X"7C",X"69",X"4D",X"2C",
		X"31",X"60",X"77",X"6E",X"43",X"2C",X"48",X"69",X"8B",X"B1",X"BA",X"9E",X"77",X"51",X"51",X"77",
		X"99",X"90",X"6E",X"80",X"A3",X"BA",X"A3",X"8B",X"A7",X"B6",X"99",X"87",X"AC",X"B1",X"90",X"69",
		X"6E",X"8B",X"AC",X"D7",X"EE",X"E0",X"B6",X"8B",X"77",X"99",X"B6",X"DB",X"E0",X"BA",X"95",X"95",
		X"B6",X"AC",X"B1",X"C4",X"BA",X"9E",X"87",X"95",X"C4",X"D2",X"B6",X"8B",X"87",X"8B",X"87",X"8B",
		X"80",X"82",X"87",X"87",X"80",X"82",X"87",X"95",X"A3",X"90",X"80",X"51",X"48",X"69",X"87",X"B1",
		X"AC",X"8B",X"6E",X"43",X"56",X"72",X"99",X"B6",X"99",X"80",X"51",X"43",X"64",X"80",X"AC",X"AC",
		X"8B",X"6E",X"43",X"4D",X"6E",X"90",X"B1",X"99",X"80",X"5B",X"31",X"22",X"3F",X"64",X"87",X"90",
		X"72",X"48",X"4D",X"6E",X"8B",X"B6",X"A3",X"82",X"60",X"3F",X"5B",X"77",X"A3",X"B1",X"90",X"77",
		X"48",X"48",X"69",X"87",X"87",X"64",X"6E",X"8B",X"80",X"60",X"77",X"95",X"BF",X"CD",X"B6",X"87",
		X"7C",X"99",X"B6",X"E5",X"DB",X"BA",X"95",X"72",X"80",X"9E",X"BA",X"A7",X"82",X"69",X"3A",X"2C",
		X"4D",X"6E",X"7C",X"56",X"5B",X"60",X"43",X"4D",X"60",X"80",X"6E",X"51",X"64",X"5B",X"3F",X"2C",
		X"48",X"77",X"7C",X"60",X"3A",X"3A",X"5B",X"7C",X"9E",X"C4",X"AC",X"90",X"69",X"4D",X"64",X"87",
		X"99",X"80",X"60",X"3A",X"14",X"14",X"3A",X"64",X"82",X"7C",X"51",X"35",X"4D",X"69",X"95",X"A7",
		X"8B",X"69",X"5B",X"69",X"51",X"51",X"69",X"69",X"51",X"56",X"6E",X"8B",X"AC",X"95",X"6E",X"5B",
		X"77",X"82",X"77",X"8B",X"90",X"80",X"64",X"3F",X"43",X"6E",X"87",X"80",X"80",X"80",X"6E",X"60",
		X"35",X"27",X"3F",X"69",X"72",X"56",X"31",X"31",X"56",X"77",X"95",X"B6",X"A7",X"87",X"69",X"4D",
		X"64",X"82",X"99",X"77",X"6E",X"87",X"AC",X"B1",X"8B",X"8B",X"AC",X"A7",X"82",X"90",X"AC",X"9E",
		X"7C",X"60",X"7C",X"9E",X"BA",X"E0",X"E9",X"C4",X"A3",X"80",X"80",X"A3",X"BF",X"E0",X"CD",X"AC",
		X"8B",X"A7",X"BA",X"A7",X"BA",X"BF",X"B1",X"90",X"87",X"AC",X"CD",X"C8",X"A3",X"80",X"8B",X"87",
		X"87",X"87",X"80",X"82",X"87",X"82",X"80",X"82",X"87",X"99",X"9E",X"8B",X"69",X"48",X"51",X"77",
		X"99",X"B6",X"A3",X"7C",X"56",X"43",X"60",X"82",X"A7",X"B1",X"90",X"69",X"48",X"48",X"6E",X"90",
		X"B1",X"A3",X"7C",X"56",X"3F",X"56",X"7C",X"A3",X"AC",X"90",X"69",X"4D",X"27",X"27",X"51",X"6E",
		X"90",X"80",X"60",X"43",X"5B",X"80",X"9E",X"B6",X"8B",X"72",X"4D",X"43",X"6E",X"87",X"AC",X"A3",
		X"80",X"60",X"3F",X"56",X"7C",X"90",X"7C",X"64",X"82",X"90",X"6E",X"69",X"87",X"A3",X"C4",X"BA",
		X"95",X"77",X"82",X"A7",X"BF",X"C4",X"A3",X"82",X"60",X"4D",X"6E",X"90",X"99",X"7C",X"51",X"35",
		X"10",X"19",X"43",X"64",X"56",X"3A",X"48",X"3A",X"2C",X"3F",X"5B",X"6E",X"48",X"48",X"4D",X"3A",
		X"1E",X"22",X"48",X"69",X"60",X"35",X"1E",X"31",X"5B",X"7C",X"9E",X"B1",X"8B",X"6E",X"48",X"43",
		X"6E",X"8B",X"87",X"64",X"3F",X"22",X"01",X"1E",X"43",X"64",X"7C",X"60",X"3A",X"31",X"51",X"77",
		X"99",X"99",X"77",X"51",X"60",X"60",X"48",X"56",X"64",X"5B",X"4D",X"5B",X"72",X"95",X"9E",X"82",
		X"60",X"5B",X"82",X"7C",X"7C",X"90",X"87",X"77",X"56",X"3F",X"51",X"77",X"87",X"80",X"82",X"7C",
		X"6E",X"4D",X"2C",X"2C",X"51",X"77",X"6E",X"4D",X"31",X"3F",X"64",X"80",X"AC",X"BF",X"9E",X"82",
		X"56",X"51",X"72",X"90",X"95",X"72",X"77",X"99",X"BF",X"A7",X"87",X"A3",X"BA",X"99",X"8B",X"AC",
		X"B1",X"95",X"69",X"6E",X"8B",X"AC",X"D7",X"EE",X"E5",X"BA",X"90",X"7C",X"90",X"B6",X"DB",X"E5",
		X"C8",X"99",X"95",X"BA",X"B6",X"B1",X"C4",X"C4",X"A7",X"87",X"99",X"BA",X"D2",X"BF",X"95",X"82",
		X"90",X"8B",X"90",X"87",X"87",X"8B",X"8B",X"82",X"87",X"8B",X"95",X"A3",X"99",X"82",X"64",X"4D",
		X"6E",X"87",X"AC",X"B6",X"90",X"77",X"51",X"56",X"77",X"95",X"B6",X"A3",X"82",X"64",X"48",X"64",
		X"82",X"A3",X"B1",X"90",X"77",X"51",X"4D",X"72",X"8B",X"B1",X"A7",X"82",X"69",X"3F",X"22",X"3F",
		X"5B",X"87",X"95",X"7C",X"56",X"4D",X"72",X"8B",X"B1",X"AC",X"87",X"69",X"48",X"5B",X"7C",X"99",
		X"B6",X"99",X"7C",X"56",X"4D",X"69",X"8B",X"90",X"69",X"6E",X"90",X"87",X"64",X"77",X"90",X"BA",
		X"C4",X"AC",X"87",X"77",X"90",X"B1",X"C4",X"B6",X"95",X"77",X"56",X"5B",X"7C",X"99",X"8B",X"64",
		X"4D",X"27",X"14",X"2C",X"51",X"64",X"3F",X"3A",X"4D",X"31",X"35",X"43",X"6E",X"60",X"3F",X"4D",
		X"4D",X"31",X"19",X"31",X"5B",X"69",X"51",X"2C",X"22",X"4D",X"6E",X"8B",X"B6",X"A3",X"87",X"60",
		X"43",X"5B",X"7C",X"90",X"7C",X"5B",X"3A",X"10",X"10",X"31",X"51",X"80",X"77",X"56",X"35",X"43",
		X"64",X"87",X"9E",X"8B",X"69",X"56",X"64",X"51",X"4D",X"60",X"69",X"51",X"51",X"69",X"8B",X"A7",
		X"9E",X"77",X"5B",X"72",X"8B",X"7C",X"8B",X"95",X"87",X"69",X"43",X"43",X"64",X"8B",X"82",X"82",
		X"82",X"77",X"69",X"43",X"2C",X"43",X"69",X"7C",X"60",X"3A",X"35",X"51",X"7C",X"99",X"BF",X"B6",
		X"90",X"72",X"51",X"64",X"8B",X"9E",X"90",X"9E",X"B6",X"D7",X"E9",X"BF",X"9E",X"7C",X"7C",X"9E",
		X"BA",X"E0",X"D2",X"A7",X"8B",X"99",X"C4",X"DB",X"BA",X"A7",X"B1",X"AC",X"B6",X"B6",X"B1",X"B1",
		X"A7",X"A7",X"B1",X"B6",X"C8",X"BF",X"A3",X"82",X"69",X"87",X"A7",X"C8",X"D7",X"B1",X"90",X"6E",
		X"6E",X"90",X"AC",X"D2",X"C4",X"95",X"80",X"8B",X"B6",X"D2",X"CD",X"C8",X"A7",X"87",X"64",X"5B",
		X"82",X"9E",X"C4",X"BA",X"90",X"77",X"56",X"69",X"90",X"A3",X"8B",X"69",X"43",X"35",X"56",X"7C",
		X"9E",X"9E",X"80",X"56",X"3A",X"43",X"69",X"8B",X"AC",X"C4",X"A7",X"87",X"69",X"56",X"7C",X"7C",
		X"77",X"7C",X"72",X"60",X"60",X"77",X"6E",X"72",X"82",X"8B",X"82",X"69",X"5B",X"64",X"56",X"3F",
		X"35",X"56",X"7C",X"7C",X"77",X"77",X"69",X"5B",X"60",X"7C",X"90",X"7C",X"56",X"35",X"22",X"4D",
		X"69",X"8B",X"90",X"6E",X"4D",X"2C",X"35",X"3A",X"3A",X"48",X"56",X"51",X"35",X"22",X"43",X"69",
		X"82",X"A7",X"AC",X"8B",X"72",X"4D",X"51",X"77",X"95",X"B1",X"9E",X"80",X"60",X"48",X"64",X"82",
		X"A3",X"B1",X"90",X"72",X"51",X"51",X"72",X"90",X"B1",X"A3",X"82",X"64",X"4D",X"60",X"82",X"95",
		X"87",X"8B",X"82",X"80",X"8B",X"99",X"9E",X"87",X"69",X"72",X"95",X"AC",X"A3",X"A7",X"A3",X"95",
		X"77",X"69",X"82",X"AC",X"B1",X"90",X"72",X"48",X"51",X"72",X"95",X"B6",X"A3",X"82",X"60",X"3A",
		X"27",X"43",X"69",X"8B",X"95",X"7C",X"51",X"51",X"72",X"90",X"BA",X"D7",X"CD",X"A3",X"80",X"60",
		X"43",X"64",X"82",X"A7",X"B6",X"8B",X"72",X"4D",X"4D",X"77",X"90",X"B6",X"A7",X"80",X"64",X"43",
		X"60",X"82",X"9E",X"BF",X"DB",X"CD",X"B1",X"82",X"87",X"A7",X"C8",X"D2",X"BA",X"9E",X"77",X"5B",
		X"72",X"8B",X"BA",X"C8",X"A7",X"82",X"7C",X"99",X"BA",X"BF",X"90",X"9E",X"99",X"99",X"A7",X"9E",
		X"9E",X"99",X"95",X"99",X"9E",X"B1",X"B6",X"A3",X"87",X"60",X"64",X"82",X"A3",X"B6",X"9E",X"82",
		X"5B",X"3F",X"5B",X"77",X"A3",X"AC",X"90",X"6E",X"64",X"82",X"A3",X"B1",X"AC",X"9E",X"80",X"5B",
		X"3A",X"51",X"6E",X"99",X"AC",X"8B",X"72",X"43",X"3F",X"60",X"80",X"82",X"64",X"43",X"22",X"31",
		X"51",X"72",X"90",X"7C",X"5B",X"3A",X"27",X"43",X"69",X"82",X"B1",X"AC",X"8B",X"6E",X"43",X"51",
		X"72",X"69",X"6E",X"69",X"5B",X"4D",X"60",X"69",X"64",X"6E",X"7C",X"82",X"72",X"51",X"56",X"5B",
		X"43",X"27",X"35",X"5B",X"72",X"6E",X"6E",X"6E",X"56",X"51",X"60",X"80",X"87",X"64",X"48",X"27",
		X"2C",X"51",X"72",X"90",X"80",X"60",X"3A",X"2C",X"35",X"31",X"3A",X"51",X"56",X"48",X"2C",X"2C",
		X"51",X"6E",X"90",X"B6",X"9E",X"82",X"5B",X"43",X"60",X"7C",X"A7",X"B1",X"90",X"77",X"48",X"4D",
		X"6E",X"8B",X"B6",X"A7",X"82",X"5B",X"43",X"5B",X"82",X"A7",X"B6",X"95",X"72",X"4D",X"4D",X"6E",
		X"95",X"87",X"8B",X"87",X"80",X"82",X"90",X"9E",X"95",X"7C",X"64",X"82",X"AC",X"AC",X"A3",X"A7",
		X"99",X"8B",X"6E",X"77",X"95",X"B6",X"A3",X"80",X"60",X"43",X"64",X"82",X"A7",X"B6",X"90",X"72",
		X"51",X"31",X"35",X"56",X"77",X"95",X"87",X"69",X"4D",X"64",X"87",X"A3",X"C8",X"D7",X"B6",X"95",
		X"77",X"4D",X"51",X"72",X"90",X"BA",X"A7",X"87",X"64",X"43",X"64",X"80",X"A7",X"B6",X"95",X"7C",
		X"4D",X"4D",X"6E",X"90",X"B6",X"D2",X"DB",X"C8",X"9E",X"82",X"95",X"BF",X"D7",X"CD",X"B6",X"8B",
		X"69",X"60",X"80",X"A7",X"C8",X"C4",X"9E",X"77",X"87",X"A7",X"C4",X"AC",X"95",X"A3",X"99",X"A3",
		X"A3",X"A3",X"A3",X"99",X"99",X"9E",X"A7",X"BA",X"B6",X"99",X"77",X"60",X"72",X"95",X"B6",X"B1",
		X"99",X"72",X"4D",X"48",X"69",X"8B",X"B1",X"AC",X"82",X"64",X"72",X"90",X"B1",X"B1",X"AC",X"95",
		X"72",X"4D",X"3F",X"60",X"82",X"A7",X"A7",X"87",X"60",X"3F",X"48",X"72",X"90",X"7C",X"60",X"35",
		X"22",X"3F",X"69",X"8B",X"90",X"72",X"48",X"2C",X"31",X"56",X"7C",X"99",X"BA",X"A3",X"7C",X"60",
		X"43",X"6E",X"72",X"69",X"72",X"64",X"56",X"51",X"69",X"69",X"69",X"77",X"82",X"80",X"64",X"51",
		X"5B",X"56",X"35",X"27",X"4D",X"72",X"72",X"6E",X"72",X"64",X"56",X"56",X"72",X"8B",X"80",X"56",
		X"31",X"1E",X"3A",X"64",X"87",X"90",X"72",X"4D",X"2C",X"31",X"35",X"35",X"43",X"56",X"51",X"35",
		X"22",X"35",X"64",X"82",X"A3",X"B6",X"8B",X"72",X"4D",X"4D",X"77",X"90",X"B6",X"A7",X"80",X"64",
		X"43",X"60",X"82",X"A3",X"B6",X"95",X"77",X"51",X"48",X"72",X"8B",X"B6",X"AC",X"82",X"69",X"48",
		X"5B",X"82",X"95",X"87",X"8B",X"82",X"82",X"87",X"99",X"9E",X"8B",X"72",X"72",X"90",X"B1",X"A7",
		X"A7",X"A3",X"99",X"80",X"69",X"82",X"A3",X"B6",X"95",X"77",X"51",X"51",X"72",X"90",X"B1",X"A7",
		X"87",X"69",X"43",X"27",X"43",X"60",X"8B",X"99",X"80",X"60",X"51",X"77",X"90",X"B6",X"DB",X"CD",
		X"AC",X"87",X"64",X"48",X"5B",X"82",X"A7",X"BA",X"9E",X"77",X"51",X"4D",X"6E",X"90",X"B6",X"AC",
		X"82",X"69",X"48",X"60",X"82",X"9E",X"BF",X"DB",X"D7",X"BA",X"95",X"8B",X"A7",X"CD",X"D7",X"BF",
		X"A3",X"80",X"64",X"72",X"90",X"B1",X"C8",X"B1",X"8B",X"7C",X"99",X"BF",X"C4",X"9E",X"9E",X"9E",
		X"99",X"A7",X"A3",X"A3",X"9E",X"99",X"99",X"A3",X"AC",X"BA",X"A7",X"90",X"6E",X"64",X"82",X"A3",
		X"B6",X"A7",X"87",X"69",X"48",X"5B",X"7C",X"99",X"B1",X"99",X"77",X"64",X"82",X"A7",X"B6",X"B1",
		X"A3",X"82",X"64",X"43",X"51",X"72",X"90",X"AC",X"95",X"77",X"51",X"43",X"60",X"82",X"8B",X"69",
		X"4D",X"27",X"2C",X"56",X"72",X"95",X"82",X"60",X"3F",X"22",X"43",X"69",X"82",X"A7",X"B1",X"90",
		X"77",X"51",X"51",X"77",X"6E",X"6E",X"6E",X"60",X"4D",X"60",X"6E",X"64",X"6E",X"80",X"82",X"77",
		X"5B",X"56",X"60",X"48",X"31",X"35",X"5B",X"77",X"72",X"72",X"6E",X"60",X"56",X"60",X"7C",X"8B",
		X"69",X"4D",X"27",X"27",X"51",X"6E",X"90",X"82",X"64",X"43",X"27",X"35",X"35",X"3A",X"4D",X"56",
		X"4D",X"2C",X"27",X"4D",X"6E",X"8B",X"AC",X"A7",X"82",X"69",X"48",X"60",X"7C",X"A3",X"B6",X"95",
		X"7C",X"4D",X"4D",X"6E",X"8B",X"B6",X"A7",X"8B",X"69",X"43",X"5B",X"7C",X"A3",X"BA",X"99",X"80",
		X"51",X"4D",X"69",X"8B",X"8B",X"8B",X"8B",X"82",X"82",X"90",X"9E",X"99",X"7C",X"69",X"7C",X"A7",
		X"B1",X"A3",X"AC",X"9E",X"90",X"72",X"72",X"95",X"B6",X"AC",X"87",X"64",X"48",X"60",X"80",X"A7",
		X"B6",X"9E",X"77",X"56",X"35",X"31",X"5B",X"77",X"99",X"90",X"69",X"51",X"5B",X"82",X"A3",X"C8",
		X"DB",X"BF",X"99",X"7C",X"56",X"51",X"72",X"90",X"B1",X"AC",X"8B",X"6E",X"4D",X"48",X"48",X"43",
		X"48",X"51",X"5B",X"51",X"4D",X"5B",X"5B",X"51",X"56",X"60",X"60",X"56",X"43",X"4D",X"60",X"82",
		X"A7",X"BA",X"A3",X"80",X"5B",X"4D",X"6E",X"90",X"B6",X"B6",X"90",X"6E",X"77",X"99",X"8B",X"95",
		X"A3",X"99",X"7C",X"6E",X"82",X"A7",X"B1",X"95",X"72",X"6E",X"77",X"77",X"7C",X"6E",X"72",X"7C",
		X"77",X"72",X"77",X"7C",X"87",X"95",X"82",X"6E",X"48",X"43",X"69",X"82",X"A7",X"A3",X"80",X"60",
		X"43",X"56",X"77",X"95",X"AC",X"90",X"77",X"51",X"48",X"69",X"87",X"B1",X"A7",X"87",X"64",X"3F",
		X"56",X"77",X"9E",X"B6",X"99",X"7C",X"56",X"31",X"27",X"48",X"72",X"95",X"90",X"72",X"4D",X"5B",
		X"7C",X"9E",X"BF",X"A3",X"87",X"5B",X"4D",X"6E",X"87",X"B6",X"B6",X"95",X"77",X"4D",X"5B",X"77",
		X"99",X"8B",X"6E",X"80",X"99",X"82",X"6E",X"87",X"AC",X"D2",X"D7",X"BA",X"8B",X"90",X"AC",X"CD",
		X"F7",X"E0",X"C4",X"99",X"7C",X"90",X"B6",X"C8",X"AC",X"8B",X"6E",X"43",X"43",X"64",X"82",X"82",
		X"60",X"6E",X"69",X"56",X"60",X"77",X"90",X"77",X"64",X"77",X"64",X"48",X"3F",X"60",X"87",X"82",
		X"64",X"48",X"4D",X"72",X"8B",X"B6",X"D2",X"B6",X"99",X"6E",X"60",X"7C",X"9E",X"A7",X"87",X"69",
		X"48",X"1E",X"2C",X"4D",X"77",X"95",X"80",X"60",X"48",X"64",X"80",X"A3",X"B1",X"95",X"72",X"6E",
		X"77",X"60",X"64",X"77",X"72",X"60",X"69",X"80",X"A3",X"B6",X"A3",X"77",X"69",X"8B",X"90",X"87",
		X"9E",X"9E",X"8B",X"69",X"4D",X"51",X"7C",X"99",X"87",X"90",X"87",X"7C",X"69",X"43",X"35",X"56",
		X"7C",X"80",X"5B",X"3A",X"3F",X"64",X"8B",X"A7",X"C4",X"AC",X"8B",X"6E",X"5B",X"77",X"99",X"A7",
		X"7C",X"80",X"99",X"BF",X"BA",X"90",X"9E",X"BF",X"AC",X"8B",X"A7",X"BA",X"A3",X"80",X"6E",X"90",
		X"B1",X"CD",X"EE",X"EE",X"C8",X"A7",X"87",X"90",X"B1",X"D2",X"EE",X"D2",X"B1",X"95",X"BA",X"C4",
		X"B1",X"C8",X"C8",X"B6",X"95",X"95",X"BF",X"D7",X"CD",X"A3",X"87",X"95",X"8B",X"90",X"8B",X"87",
		X"8B",X"90",X"87",X"87",X"8B",X"95",X"A7",X"A3",X"8B",X"6E",X"51",X"60",X"82",X"AC",X"BF",X"A3",
		X"80",X"56",X"4D",X"6E",X"90",X"B6",X"B1",X"90",X"69",X"4D",X"56",X"7C",X"A3",X"BA",X"A3",X"7C",
		X"56",X"48",X"64",X"8B",X"B1",X"B1",X"90",X"69",X"4D",X"27",X"35",X"60",X"7C",X"99",X"82",X"60",
		X"4D",X"64",X"87",X"AC",X"B6",X"95",X"72",X"4D",X"51",X"72",X"99",X"B6",X"A7",X"82",X"5B",X"48",
		X"5B",X"87",X"99",X"77",X"69",X"8B",X"90",X"6E",X"6E",X"90",X"B1",X"C8",X"BA",X"90",X"77",X"82",
		X"AC",X"C8",X"BF",X"A7",X"80",X"5B",X"51",X"72",X"99",X"95",X"77",X"56",X"2C",X"14",X"1E",X"4D",
		X"69",X"4D",X"3A",X"4D",X"35",X"31",X"43",X"64",X"69",X"48",X"4D",X"4D",X"3A",X"1E",X"2C",X"56",
		X"6E",X"5B",X"31",X"22",X"3A",X"69",X"82",X"A7",X"B1",X"87",X"6E",X"48",X"51",X"77",X"90",X"87",
		X"60",X"3F",X"1E",X"06",X"2C",X"4D",X"72",X"80",X"5B",X"3A",X"35",X"5B",X"82",X"9E",X"95",X"72",
		X"51",X"64",X"5B",X"4D",X"5B",X"69",X"5B",X"51",X"64",X"7C",X"9E",X"9E",X"80",X"5B",X"69",X"8B",
		X"7C",X"82",X"95",X"87",X"77",X"51",X"3F",X"5B",X"82",X"87",X"80",X"82",X"7C",X"6E",X"48",X"2C",
		X"31",X"60",X"7C",X"69",X"48",X"31",X"4D",X"6E",X"8B",X"B6",X"BA",X"99",X"7C",X"51",X"5B",X"7C",
		X"99",X"90",X"72",X"80",X"A7",X"BF",X"A3",X"8B",X"AC",X"BA",X"95",X"8B",X"B6",X"B1",X"90",X"72",
		X"72",X"95",X"B1",X"DB",X"F7",X"DB",X"BA",X"90",X"80",X"99",X"B6",X"E5",X"E5",X"C4",X"9E",X"99",
		X"C4",X"B6",X"B6",X"C8",X"BF",X"A7",X"8B",X"9E",X"C4",X"D7",X"BA",X"8B",X"87",X"90",X"8B",X"90",
		X"87",X"87",X"8B",X"8B",X"82",X"87",X"8B",X"99",X"A7",X"99",X"80",X"60",X"4D",X"72",X"90",X"B1",
		X"B1",X"8B",X"72",X"4D",X"60",X"80",X"9E",X"B6",X"9E",X"80",X"5B",X"4D",X"6E",X"87",X"AC",X"B1",
		X"8B",X"72",X"4D",X"56",X"77",X"95",X"B1",X"9E",X"7C",X"60",X"35",X"27",X"48",X"64",X"90",X"90",
		X"77",X"51",X"51",X"77",X"95",X"B6",X"A3",X"82",X"64",X"48",X"64",X"82",X"A3",X"B1",X"90",X"77",
		X"51",X"51",X"6E",X"90",X"8B",X"64",X"77",X"95",X"80",X"64",X"80",X"99",X"BF",X"C4",X"A7",X"82",
		X"7C",X"95",X"B6",X"C4",X"AC",X"90",X"72",X"51",X"60",X"82",X"9E",X"82",X"60",X"43",X"1E",X"14",
		X"31",X"5B",X"64",X"3A",X"43",X"48",X"31",X"3A",X"4D",X"72",X"56",X"3F",X"51",X"48",X"27",X"19",
		X"3A",X"60",X"69",X"48",X"27",X"27",X"51",X"72",X"90",X"B1",X"9E",X"80",X"60",X"48",X"60",X"82",
		X"95",X"72",X"51",X"35",X"14",X"14",X"35",X"56",X"7C",X"72",X"51",X"31",X"48",X"6E",X"8B",X"A3",
		X"87",X"60",X"5B",X"69",X"4D",X"51",X"64",X"69",X"4D",X"5B",X"69",X"8B",X"AC",X"95",X"77",X"5B",
		X"7C",X"87",X"77",X"90",X"90",X"82",X"69",X"3F",X"48",X"69",X"87",X"82",X"82",X"82",X"72",X"64",
		X"3A",X"31",X"48",X"72",X"7C",X"56",X"35",X"35",X"5B",X"82",X"9E",X"C4",X"AC",X"87",X"6E",X"4D",
		X"6E",X"90",X"A3",X"80",X"77",X"90",X"B6",X"BA",X"90",X"99",X"BA",X"AC",X"87",X"9E",X"BA",X"A3",
		X"7C",X"6E",X"80",X"A7",X"C8",X"E9",X"F3",X"C8",X"A7",X"82",X"87",X"B1",X"C8",X"EE",X"D7",X"AC",
		X"95",X"AC",X"BF",X"B1",X"C4",X"C8",X"B6",X"95",X"90",X"B1",X"D7",X"CD",X"A7",X"8B",X"90",X"8B",
		X"90",X"8B",X"87",X"8B",X"90",X"87",X"82",X"8B",X"90",X"A7",X"A3",X"90",X"77",X"4D",X"60",X"7C",
		X"A3",X"BF",X"A3",X"87",X"5B",X"4D",X"6E",X"87",X"B6",X"B6",X"95",X"77",X"48",X"56",X"77",X"99",
		X"BA",X"A3",X"87",X"60",X"48",X"64",X"80",X"AC",X"B1",X"95",X"77",X"4D",X"2C",X"31",X"56",X"7C",
		X"99",X"8B",X"64",X"48",X"64",X"80",X"A7",X"BA",X"99",X"7C",X"4D",X"51",X"6E",X"8B",X"BA",X"A7",
		X"8B",X"64",X"43",X"5B",X"7C",X"95",X"7C",X"69",X"82",X"90",X"72",X"69",X"87",X"B1",X"C8",X"BF",
		X"99",X"72",X"82",X"A3",X"C4",X"BF",X"A7",X"87",X"60",X"51",X"6E",X"95",X"99",X"77",X"56",X"31",
		X"14",X"1E",X"48",X"69",X"51",X"35",X"48",X"3A",X"31",X"3F",X"64",X"6E",X"48",X"48",X"4D",X"3F",
		X"1E",X"27",X"56",X"6E",X"64",X"3A",X"22",X"3A",X"60",X"82",X"A7",X"B1",X"95",X"6E",X"4D",X"4D",
		X"6E",X"95",X"87",X"69",X"48",X"1E",X"0B",X"1E",X"48",X"72",X"80",X"69",X"3A",X"35",X"5B",X"77",
		X"A3",X"99",X"7C",X"5B",X"64",X"60",X"4D",X"5B",X"6E",X"60",X"51",X"64",X"7C",X"9E",X"A7",X"82",
		X"64",X"64",X"82",X"80",X"80",X"95",X"8B",X"77",X"56",X"3F",X"56",X"80",X"8B",X"80",X"87",X"7C",
		X"72",X"51",X"2C",X"35",X"56",X"77",X"6E",X"4D",X"31",X"48",X"6E",X"87",X"AC",X"BF",X"9E",X"80",
		X"60",X"5B",X"7C",X"99",X"99",X"95",X"AC",X"C4",X"E5",X"CD",X"AC",X"8B",X"77",X"90",X"AC",X"D2",
		X"DB",X"BA",X"95",X"90",X"B6",X"D7",X"CD",X"A7",X"B6",X"AC",X"B1",X"B6",X"B1",X"B6",X"AC",X"A7",
		X"AC",X"B1",X"BF",X"C4",X"B1",X"95",X"72",X"7C",X"99",X"BA",X"D7",X"BF",X"9E",X"80",X"69",X"82",
		X"9E",X"C4",X"CD",X"AC",X"87",X"82",X"AC",X"C8",X"D2",X"CD",X"B6",X"95",X"6E",X"56",X"77",X"90",
		X"BA",X"C4",X"A3",X"82",X"56",X"60",X"80",X"9E",X"95",X"72",X"56",X"35",X"4D",X"6E",X"90",X"A3",
		X"87",X"69",X"43",X"3A",X"60",X"7C",X"9E",X"C4",X"B6",X"95",X"72",X"51",X"69",X"82",X"77",X"7C",
		X"77",X"64",X"5B",X"72",X"72",X"6E",X"7C",X"87",X"8B",X"77",X"56",X"64",X"64",X"43",X"31",X"43",
		X"6E",X"7C",X"72",X"77",X"72",X"5B",X"5B",X"6E",X"87",X"87",X"64",X"48",X"27",X"3A",X"5B",X"80",
		X"95",X"7C",X"60",X"3A",X"31",X"3A",X"35",X"43",X"56",X"56",X"43",X"2C",X"31",X"5B",X"77",X"9E",
		X"B6",X"99",X"80",X"51",X"48",X"69",X"82",X"B1",X"AC",X"8B",X"6E",X"43",X"56",X"72",X"99",X"B6",
		X"9E",X"82",X"56",X"43",X"64",X"80",X"AC",X"B1",X"90",X"72",X"48",X"51",X"72",X"90",X"87",X"8B",
		X"87",X"80",X"82",X"90",X"9E",X"90",X"72",X"69",X"82",X"AC",X"A7",X"A3",X"A7",X"95",X"87",X"64",
		X"77",X"9E",X"B6",X"9E",X"7C",X"56",X"43",X"64",X"87",X"AC",X"B1",X"90",X"69",X"4D",X"27",X"35",
		X"5B",X"7C",X"99",X"82",X"5B",X"48",X"69",X"8B",X"A7",X"CD",X"CD",X"AC",X"8B",X"6E",X"43",X"56",
		X"72",X"99",X"B6",X"9E",X"80",X"56",X"43",X"64",X"80",X"AC",X"B1",X"90",X"72",X"43",X"51",X"72",
		X"95",X"BA",X"D7",X"D7",X"BA",X"95",X"82",X"95",X"C4",X"D2",X"C8",X"A7",X"80",X"60",X"64",X"82",
		X"AC",X"C8",X"BA",X"90",X"72",X"8B",X"AC",X"C4",X"9E",X"95",X"9E",X"95",X"A3",X"9E",X"9E",X"9E",
		X"95",X"95",X"99",X"A7",X"B6",X"AC",X"90",X"6E",X"5B",X"72",X"99",X"B1",X"AC",X"8B",X"69",X"43",
		X"48",X"6E",X"95",X"AC",X"A3",X"7C",X"60",X"77",X"95",X"B1",X"AC",X"A7",X"8B",X"64",X"43",X"3F",
		X"64",X"87",X"A7",X"9E",X"7C",X"51",X"3A",X"4D",X"77",X"8B",X"72",X"56",X"27",X"22",X"43",X"64",
		X"90",X"87",X"69",X"48",X"22",X"35",X"56",X"7C",X"9E",X"B6",X"9E",X"77",X"51",X"43",X"69",X"6E",
		X"69",X"6E",X"60",X"4D",X"56",X"69",X"64",X"69",X"77",X"82",X"7C",X"5B",X"4D",X"5B",X"4D",X"2C",
		X"27",X"48",X"77",X"6E",X"6E",X"6E",X"60",X"51",X"56",X"77",X"8B",X"72",X"56",X"2C",X"1E",X"3F",
		X"60",X"8B",X"8B",X"69",X"43",X"27",X"31",X"35",X"35",X"48",X"56",X"4D",X"31",X"22",X"3F",X"69",
		X"87",X"A7",X"AC",X"82",X"69",X"43",X"51",X"7C",X"95",X"B6",X"99",X"7C",X"5B",X"43",X"64",X"82",
		X"A7",X"B1",X"8B",X"6E",X"48",X"4D",X"77",X"90",X"B6",X"A3",X"80",X"60",X"43",X"60",X"87",X"90",
		X"87",X"8B",X"80",X"80",X"87",X"9E",X"99",X"87",X"6E",X"77",X"99",X"B1",X"A7",X"A7",X"9E",X"95",
		X"77",X"69",X"87",X"A7",X"B1",X"8B",X"72",X"4D",X"56",X"77",X"95",X"B1",X"A3",X"80",X"64",X"3A",
		X"27",X"48",X"69",X"90",X"95",X"77",X"56",X"56",X"7C",X"95",X"BA",X"DB",X"C4",X"A3",X"80",X"5B",
		X"48",X"64",X"87",X"AC",X"B6",X"95",X"72",X"4D",X"51",X"72",X"99",X"B6",X"A7",X"82",X"60",X"48",
		X"60",X"82",X"A7",X"C4",X"DB",X"CD",X"B1",X"8B",X"87",X"B1",X"CD",X"D7",X"BF",X"99",X"7C",X"5B",
		X"77",X"95",X"BA",X"CD",X"A7",X"82",X"7C",X"99",X"BF",X"BF",X"95",X"9E",X"9E",X"9E",X"A7",X"A3",
		X"A3",X"9E",X"95",X"99",X"A3",X"B1",X"BA",X"A3",X"87",X"64",X"64",X"8B",X"A7",X"B6",X"A3",X"80",
		X"60",X"43",X"60",X"80",X"A3",X"AC",X"90",X"6E",X"64",X"8B",X"A7",X"B1",X"AC",X"99",X"7C",X"5B",
		X"3F",X"56",X"77",X"95",X"AC",X"8B",X"72",X"48",X"43",X"64",X"87",X"87",X"60",X"43",X"1E",X"31",
		X"5B",X"77",X"95",X"7C",X"5B",X"35",X"27",X"48",X"6E",X"87",X"AC",X"AC",X"87",X"6E",X"48",X"56",
		X"77",X"69",X"6E",X"69",X"5B",X"4D",X"64",X"69",X"64",X"6E",X"80",X"82",X"72",X"56",X"56",X"5B",
		X"43",X"2C",X"3A",X"64",X"77",X"6E",X"72",X"6E",X"5B",X"56",X"64",X"82",X"87",X"60",X"43",X"22",
		X"2C",X"56",X"72",X"95",X"7C",X"5B",X"3A",X"27",X"35",X"35",X"3F",X"4D",X"56",X"48",X"27",X"2C",
		X"56",X"72",X"95",X"B1",X"9E",X"80",X"60",X"48",X"64",X"82",X"A3",X"B1",X"90",X"72",X"4D",X"51",
		X"72",X"90",X"B1",X"A3",X"82",X"64",X"48",X"60",X"80",X"A3",X"B6",X"95",X"77",X"51",X"51",X"6E",
		X"90",X"90",X"8B",X"8B",X"80",X"82",X"95",X"9E",X"99",X"77",X"69",X"82",X"A7",X"AC",X"A7",X"AC",
		X"9E",X"8B",X"6E",X"72",X"95",X"BA",X"A3",X"87",X"60",X"48",X"64",X"80",X"AC",X"B6",X"95",X"6E",
		X"51",X"2C",X"35",X"60",X"7C",X"9E",X"87",X"64",X"4D",X"64",X"8B",X"AC",X"CD",X"DB",X"B6",X"90",
		X"77",X"51",X"56",X"77",X"95",X"B6",X"A7",X"82",X"64",X"4D",X"64",X"82",X"A7",X"B6",X"95",X"77",
		X"51",X"51",X"72",X"90",X"B1",X"DB",X"DB",X"C8",X"9E",X"82",X"99",X"BA",X"D7",X"CD",X"B1",X"90",
		X"64",X"64",X"82",X"A3",X"CD",X"BF",X"9E",X"7C",X"8B",X"AC",X"C8",X"A7",X"95",X"A3",X"95",X"A7",
		X"A3",X"A3",X"A3",X"99",X"99",X"9E",X"A7",X"BA",X"B1",X"9E",X"77",X"5B",X"77",X"95",X"B1",X"B1",
		X"95",X"77",X"48",X"4D",X"69",X"8B",X"B1",X"A3",X"82",X"69",X"77",X"95",X"B1",X"B1",X"AC",X"90",
		X"72",X"48",X"3F",X"64",X"80",X"AC",X"A3",X"82",X"60",X"3A",X"51",X"72",X"8B",X"77",X"56",X"35",
		X"22",X"43",X"64",X"87",X"8B",X"6E",X"4D",X"2C",X"31",X"56",X"77",X"99",X"BA",X"9E",X"82",X"5B",
		X"43",X"69",X"72",X"6E",X"6E",X"69",X"56",X"56",X"69",X"69",X"69",X"77",X"82",X"82",X"60",X"4D",
		X"60",X"56",X"35",X"27",X"48",X"6E",X"72",X"6E",X"72",X"64",X"56",X"56",X"72",X"8B",X"77",X"5B",
		X"31",X"1E",X"43",X"60",X"8B",X"8B",X"72",X"51",X"27",X"35",X"35",X"35",X"48",X"56",X"56",X"35",
		X"22",X"3F",X"60",X"82",X"A7",X"B1",X"90",X"6E",X"4D",X"4D",X"72",X"95",X"B6",X"A7",X"82",X"5B",
		X"48",X"5B",X"82",X"A7",X"B6",X"99",X"72",X"51",X"4D",X"6E",X"95",X"B6",X"AC",X"87",X"60",X"48",
		X"56",X"82",X"95",X"87",X"90",X"82",X"82",X"87",X"99",X"9E",X"8B",X"6E",X"72",X"99",X"B1",X"A7",
		X"A7",X"A3",X"95",X"80",X"6E",X"82",X"A7",X"B6",X"90",X"77",X"4D",X"4D",X"77",X"90",X"B6",X"A7",
		X"82",X"64",X"43",X"2C",X"43",X"64",X"87",X"95",X"7C",X"56",X"51",X"7C",X"95",X"B6",X"D7",X"CD",
		X"A7",X"8B",X"64",X"48",X"64",X"80",X"A7",X"BA",X"99",X"7C",X"51",X"48",X"48",X"48",X"4D",X"4D",
		X"4D",X"51",X"51",X"51",X"51",X"56",X"56",X"56",X"56",X"5B",X"5B",X"5B",X"5B",X"5B",X"60",X"60",
		X"60",X"60",X"60",X"64",X"64",X"64",X"64",X"64",X"64",X"69",X"69",X"69",X"69",X"69",X"69",X"6E",
		X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"77",
		X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"82",X"82",X"87",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"7C",X"7C",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"7C",X"80",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"80",
		X"7C",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"7C",X"80",
		X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"80",X"80",X"7C",X"7C",X"80",
		X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"7C",X"7C",
		X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"80",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"80",X"80",
		X"80",X"80",X"7C",X"80",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"7C",X"72",X"77",X"7C",X"7C",X"7C",X"77",X"72",
		X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"80",X"77",X"77",X"7C",X"7C",X"7C",X"82",X"80",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",
		X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",
		X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",
		X"80",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",
		X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"82",X"80",X"77",
		X"80",X"82",X"80",X"77",X"80",X"82",X"7C",X"77",X"82",X"82",X"77",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",
		X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"72",X"77",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",
		X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"80",
		X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"72",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"7C",
		X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"7C",X"7C",
		X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",
		X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",
		X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"80",X"82",
		X"80",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"77",X"80",
		X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",
		X"7C",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",
		X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"72",
		X"77",X"80",X"87",X"7C",X"77",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",
		X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"82",X"80",X"77",X"7C",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"72",X"7C",X"7C",X"7C",X"7C",X"77",
		X"77",X"7C",X"7C",X"7C",X"7C",X"77",X"7C",X"80",X"77",X"77",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",
		X"80",X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"7C",X"82",X"82",X"80",X"7C",X"7C",X"7C",
		X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"82",
		X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"8B",X"82",X"8B",X"8B",X"8B",X"90",X"90",X"90",X"95",
		X"95",X"95",X"95",X"95",X"90",X"95",X"99",X"95",X"90",X"87",X"8B",X"87",X"80",X"7C",X"80",X"7C",
		X"72",X"72",X"72",X"6E",X"64",X"69",X"64",X"60",X"51",X"43",X"4D",X"48",X"51",X"56",X"51",X"51",
		X"51",X"51",X"56",X"64",X"60",X"64",X"69",X"69",X"6E",X"72",X"72",X"72",X"80",X"80",X"7C",X"82",
		X"8B",X"8B",X"87",X"90",X"99",X"95",X"95",X"99",X"99",X"90",X"95",X"99",X"95",X"8B",X"87",X"8B",
		X"82",X"7C",X"7C",X"80",X"77",X"77",X"77",X"6E",X"72",X"6E",X"69",X"6E",X"77",X"7C",X"72",X"6E",
		X"7C",X"7C",X"7C",X"80",X"87",X"87",X"7C",X"80",X"87",X"82",X"87",X"8B",X"87",X"82",X"82",X"80",
		X"7C",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"7C",X"80",X"82",X"82",X"82",X"80",X"87",
		X"87",X"87",X"87",X"87",X"87",X"82",X"80",X"87",X"82",X"87",X"8B",X"87",X"82",X"7C",X"82",X"87",
		X"80",X"7C",X"80",X"7C",X"77",X"77",X"7C",X"77",X"77",X"80",X"80",X"77",X"7C",X"77",X"72",X"77",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"72",X"72",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"72",
		X"77",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",
		X"80",X"7C",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",X"80",X"80",X"80",X"80",X"77",X"7C",
		X"77",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"7C",
		X"72",X"77",X"7C",X"7C",X"7C",X"7C",X"80",X"77",X"77",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",
		X"77",X"80",X"7C",X"77",X"77",X"77",X"77",X"77",X"7C",X"82",X"87",X"7C",X"7C",X"80",X"77",X"77",
		X"80",X"87",X"82",X"82",X"80",X"77",X"77",X"7C",X"87",X"95",X"7C",X"80",X"80",X"7C",X"82",X"80",
		X"82",X"87",X"87",X"80",X"77",X"80",X"82",X"80",X"87",X"87",X"82",X"7C",X"7C",X"7C",X"7C",X"80",
		X"80",X"82",X"80",X"7C",X"7C",X"77",X"72",X"77",X"80",X"82",X"7C",X"7C",X"7C",X"72",X"77",X"7C",
		X"82",X"80",X"77",X"7C",X"7C",X"72",X"77",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",
		X"80",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"72",X"7C",X"7C",X"7C",X"7C",X"77",X"77",
		X"77",X"77",X"80",X"7C",X"80",X"7C",X"80",X"7C",X"77",X"7C",X"80",X"7C",X"80",X"77",X"77",X"7C",
		X"82",X"82",X"7C",X"80",X"87",X"82",X"7C",X"80",X"87",X"82",X"82",X"82",X"82",X"80",X"7C",X"80",
		X"82",X"7C",X"7C",X"82",X"80",X"82",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"82",
		X"7C",X"7C",X"82",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"80",
		X"72",X"72",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"72",X"77",X"80",X"77",X"72",X"7C",X"80",X"7C",
		X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"7C",X"77",X"77",X"80",X"7C",X"80",X"82",X"80",X"77",X"72",
		X"7C",X"80",X"7C",X"82",X"82",X"7C",X"80",X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",
		X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"82",X"80",X"7C",X"80",X"82",X"80",
		X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"82",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"80",
		X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"77",
		X"72",X"7C",X"80",X"7C",X"80",X"82",X"80",X"77",X"77",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",
		X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"7C",X"7C",X"82",X"80",X"7C",
		X"7C",X"7C",X"72",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",
		X"7C",X"80",X"7C",X"80",X"82",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"82",X"7C",X"7C",X"82",
		X"80",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"80",X"80",X"80",X"7C",X"7C",X"80",
		X"80",X"7C",X"7C",X"80",X"80",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",
		X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",
		X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",
		X"80",X"80",X"7C",X"7C",X"80",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"7C",X"7C",X"80",X"82",X"7C",
		X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",
		X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",
		X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"77",X"80",X"82",X"7C",X"7C",X"80",
		X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"77",X"7C",X"82",X"7C",
		X"77",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"77",X"7C",X"82",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",
		X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",
		X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",
		X"82",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",
		X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",
		X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",
		X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"7C",
		X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",
		X"82",X"82",X"7C",X"7C",X"80",X"87",X"87",X"7C",X"80",X"87",X"82",X"7C",X"82",X"87",X"82",X"77",
		X"69",X"7C",X"95",X"B1",X"D7",X"D7",X"B1",X"95",X"72",X"7C",X"99",X"BF",X"DB",X"BF",X"9E",X"82",
		X"A7",X"AC",X"9E",X"B6",X"B6",X"A3",X"87",X"87",X"A7",X"C8",X"BA",X"8B",X"7C",X"82",X"82",X"82",
		X"80",X"7C",X"82",X"82",X"7C",X"7C",X"82",X"87",X"99",X"95",X"80",X"64",X"43",X"5B",X"80",X"99",
		X"B6",X"90",X"72",X"51",X"43",X"6E",X"87",X"AC",X"A7",X"82",X"64",X"43",X"51",X"7C",X"95",X"B6",
		X"95",X"77",X"51",X"3F",X"69",X"82",X"A7",X"AC",X"82",X"69",X"48",X"27",X"31",X"56",X"77",X"90",
		X"80",X"5B",X"43",X"64",X"82",X"A7",X"B1",X"8B",X"6E",X"48",X"4D",X"77",X"90",X"B6",X"9E",X"7C",
		X"60",X"43",X"60",X"82",X"95",X"77",X"69",X"87",X"90",X"6E",X"6E",X"8B",X"AC",X"CD",X"BF",X"99",
		X"7C",X"90",X"B6",X"D2",X"E9",X"BF",X"A3",X"7C",X"72",X"95",X"B6",X"B6",X"90",X"6E",X"4D",X"2C",
		X"3F",X"69",X"80",X"69",X"51",X"64",X"51",X"48",X"5B",X"7C",X"80",X"5B",X"60",X"60",X"4D",X"31",
		X"3F",X"64",X"80",X"6E",X"3F",X"31",X"48",X"77",X"90",X"B6",X"BF",X"95",X"7C",X"56",X"5B",X"80",
		X"99",X"90",X"6E",X"48",X"27",X"10",X"31",X"51",X"77",X"80",X"64",X"3F",X"3F",X"69",X"82",X"A7",
		X"99",X"72",X"5B",X"69",X"60",X"4D",X"60",X"6E",X"5B",X"51",X"64",X"7C",X"AC",X"A3",X"82",X"64",
		X"6E",X"8B",X"7C",X"82",X"95",X"87",X"7C",X"4D",X"3F",X"5B",X"80",X"82",X"80",X"82",X"77",X"69",
		X"48",X"27",X"35",X"64",X"77",X"6E",X"3F",X"2C",X"48",X"69",X"90",X"B6",X"BA",X"99",X"72",X"51",
		X"56",X"7C",X"9E",X"8B",X"6E",X"80",X"A7",X"BA",X"A3",X"8B",X"A7",X"B6",X"95",X"8B",X"AC",X"B1",
		X"8B",X"64",X"72",X"90",X"B1",X"DB",X"EE",X"DB",X"B1",X"8B",X"7C",X"95",X"BA",X"DB",X"E0",X"BF",
		X"95",X"95",X"BF",X"B1",X"B6",X"C4",X"BF",X"9E",X"87",X"99",X"BF",X"CD",X"B6",X"8B",X"82",X"8B",
		X"87",X"8B",X"82",X"82",X"87",X"87",X"80",X"82",X"87",X"95",X"A3",X"95",X"80",X"5B",X"4D",X"6E",
		X"87",X"AC",X"AC",X"8B",X"6E",X"4D",X"56",X"77",X"95",X"B1",X"99",X"7C",X"5B",X"48",X"64",X"82",
		X"A7",X"AC",X"87",X"6E",X"48",X"51",X"72",X"90",X"AC",X"9E",X"7C",X"60",X"35",X"22",X"43",X"60",
		X"8B",X"8B",X"72",X"4D",X"4D",X"72",X"90",X"B6",X"9E",X"82",X"5B",X"43",X"60",X"7C",X"A7",X"B1",
		X"90",X"72",X"43",X"4D",X"69",X"8B",X"82",X"64",X"72",X"90",X"7C",X"60",X"77",X"99",X"BF",X"BF",
		X"A3",X"77",X"77",X"90",X"B1",X"C4",X"AC",X"90",X"69",X"48",X"5B",X"80",X"95",X"82",X"60",X"43",
		X"14",X"10",X"31",X"51",X"5B",X"35",X"3F",X"43",X"2C",X"35",X"48",X"69",X"51",X"3F",X"4D",X"43",
		X"27",X"19",X"35",X"64",X"69",X"48",X"27",X"27",X"4D",X"6E",X"90",X"B1",X"99",X"80",X"56",X"3F",
		X"5B",X"80",X"8B",X"72",X"51",X"31",X"06",X"10",X"31",X"56",X"80",X"6E",X"4D",X"31",X"48",X"69",
		X"8B",X"9E",X"82",X"60",X"56",X"64",X"4D",X"4D",X"60",X"64",X"4D",X"56",X"69",X"90",X"A7",X"95",
		X"6E",X"56",X"77",X"87",X"7C",X"8B",X"90",X"82",X"60",X"3F",X"43",X"69",X"8B",X"80",X"82",X"80",
		X"72",X"60",X"3A",X"2C",X"43",X"6E",X"7C",X"56",X"35",X"35",X"56",X"80",X"99",X"BF",X"AC",X"87",
		X"6E",X"4D",X"69",X"8B",X"9E",X"80",X"77",X"90",X"B6",X"BA",X"90",X"95",X"B6",X"AC",X"87",X"99",
		X"B6",X"A3",X"7C",X"69",X"82",X"A7",X"C4",X"E5",X"EE",X"C8",X"A7",X"82",X"87",X"AC",X"C8",X"E9",
		X"D2",X"B1",X"90",X"B1",X"BF",X"AC",X"BF",X"C4",X"B6",X"95",X"8B",X"B6",X"D2",X"CD",X"A3",X"82",
		X"90",X"8B",X"8B",X"8B",X"82",X"8B",X"8B",X"87",X"82",X"8B",X"90",X"A3",X"A3",X"90",X"6E",X"4D",
		X"5B",X"80",X"A3",X"BA",X"A7",X"80",X"5B",X"4D",X"69",X"8B",X"B1",X"B6",X"90",X"6E",X"4D",X"51",
		X"77",X"9E",X"B6",X"A7",X"80",X"5B",X"48",X"60",X"82",X"AC",X"B1",X"95",X"6E",X"51",X"2C",X"31",
		X"5B",X"77",X"99",X"87",X"60",X"48",X"60",X"82",X"A7",X"B6",X"99",X"77",X"51",X"4D",X"6E",X"95",
		X"B6",X"AC",X"87",X"60",X"48",X"56",X"80",X"99",X"7C",X"64",X"87",X"95",X"72",X"69",X"8B",X"AC",
		X"C4",X"BA",X"90",X"77",X"80",X"A7",X"C4",X"BF",X"A7",X"82",X"5B",X"51",X"69",X"95",X"99",X"7C",
		X"5B",X"31",X"14",X"19",X"43",X"69",X"51",X"35",X"48",X"3A",X"31",X"3F",X"60",X"6E",X"48",X"48",
		X"51",X"3F",X"1E",X"22",X"51",X"6E",X"64",X"3A",X"22",X"3A",X"5B",X"80",X"A7",X"B1",X"8B",X"72",
		X"4D",X"4D",X"77",X"90",X"8B",X"64",X"43",X"22",X"06",X"27",X"48",X"6E",X"80",X"60",X"3A",X"35",
		X"56",X"80",X"9E",X"99",X"77",X"56",X"64",X"60",X"4D",X"5B",X"69",X"60",X"51",X"64",X"77",X"9E",
		X"A3",X"87",X"64",X"64",X"8B",X"80",X"80",X"95",X"8B",X"7C",X"56",X"43",X"56",X"80",X"8B",X"80",
		X"87",X"7C",X"72",X"4D",X"2C",X"31",X"5B",X"7C",X"6E",X"4D",X"31",X"48",X"6E",X"87",X"B1",X"BF",
		X"9E",X"82",X"56",X"5B",X"77",X"99",X"95",X"72",X"80",X"A3",X"C4",X"A7",X"8B",X"A7",X"BF",X"9E",
		X"8B",X"B1",X"B6",X"95",X"77",X"72",X"95",X"B1",X"D7",X"F7",X"E0",X"BF",X"99",X"80",X"99",X"B1",
		X"E0",X"E9",X"C8",X"A7",X"99",X"BF",X"B6",X"B6",X"CD",X"C4",X"AC",X"90",X"9E",X"C4",X"DB",X"BF",
		X"95",X"87",X"95",X"8B",X"90",X"87",X"87",X"90",X"8B",X"87",X"87",X"90",X"95",X"A7",X"9E",X"82",
		X"64",X"4D",X"72",X"8B",X"B1",X"BA",X"90",X"77",X"51",X"56",X"80",X"99",X"BA",X"A7",X"82",X"64",
		X"48",X"69",X"87",X"A7",X"BA",X"90",X"77",X"51",X"4D",X"77",X"90",X"B1",X"A7",X"82",X"69",X"3F",
		X"27",X"48",X"64",X"90",X"95",X"7C",X"5B",X"51",X"77",X"90",X"B6",X"AC",X"87",X"69",X"4D",X"60",
		X"80",X"9E",X"B6",X"99",X"7C",X"56",X"51",X"6E",X"90",X"90",X"69",X"72",X"95",X"87",X"64",X"7C",
		X"95",X"BF",X"C8",X"AC",X"87",X"7C",X"95",X"B6",X"C8",X"B6",X"95",X"77",X"56",X"60",X"80",X"9E",
		X"8B",X"64",X"4D",X"27",X"14",X"31",X"56",X"69",X"3F",X"3F",X"4D",X"31",X"3A",X"48",X"6E",X"60",
		X"3F",X"51",X"4D",X"2C",X"19",X"35",X"5B",X"6E",X"51",X"2C",X"27",X"51",X"6E",X"8B",X"B1",X"A3",
		X"82",X"64",X"48",X"5B",X"80",X"95",X"7C",X"56",X"3A",X"19",X"10",X"35",X"51",X"7C",X"77",X"56",
		X"31",X"43",X"69",X"87",X"A7",X"8B",X"64",X"56",X"69",X"51",X"4D",X"64",X"69",X"51",X"56",X"69",
		X"87",X"AC",X"99",X"7C",X"60",X"77",X"8B",X"7C",X"8B",X"95",X"87",X"72",X"43",X"43",X"64",X"87",
		X"82",X"82",X"82",X"77",X"64",X"43",X"27",X"43",X"6E",X"7C",X"64",X"3A",X"35",X"56",X"77",X"9E",
		X"BF",X"B6",X"95",X"6E",X"51",X"60",X"8B",X"A3",X"90",X"9E",X"B6",X"DB",X"E5",X"BA",X"9E",X"7C",
		X"7C",X"A3",X"BF",X"E0",X"CD",X"A3",X"8B",X"9E",X"C8",X"DB",X"B6",X"A7",X"B1",X"AC",X"BA",X"B6",
		X"B6",X"B1",X"A7",X"AC",X"B1",X"BA",X"CD",X"BF",X"A3",X"82",X"6E",X"8B",X"AC",X"CD",X"D7",X"AC",
		X"90",X"69",X"72",X"95",X"B1",X"D2",X"BF",X"95",X"80",X"90",X"BA",X"D2",X"CD",X"C8",X"A3",X"87",
		X"64",X"60",X"87",X"A3",X"C8",X"B6",X"90",X"72",X"56",X"6E",X"90",X"A3",X"8B",X"64",X"3F",X"35",
		X"5B",X"80",X"9E",X"9E",X"7C",X"56",X"3A",X"43",X"6E",X"8B",X"AC",X"C8",X"A7",X"82",X"64",X"51",
		X"80",X"7C",X"77",X"7C",X"6E",X"5B",X"60",X"72",X"6E",X"72",X"80",X"8B",X"82",X"69",X"5B",X"64",
		X"56",X"3A",X"31",X"5B",X"7C",X"77",X"72",X"77",X"69",X"5B",X"60",X"7C",X"90",X"80",X"56",X"31",
		X"27",X"43",X"6E",X"90",X"90",X"72",X"4D",X"2C",X"35",X"3A",X"3A",X"4D",X"5B",X"51",X"35",X"27",
		X"3F",X"69",X"87",X"AC",X"B1",X"87",X"6E",X"48",X"51",X"7C",X"95",X"B6",X"9E",X"7C",X"60",X"43",
		X"64",X"82",X"A7",X"B6",X"8B",X"72",X"4D",X"51",X"77",X"90",X"B1",X"9E",X"82",X"60",X"48",X"60",
		X"87",X"90",X"87",X"8B",X"80",X"80",X"8B",X"99",X"99",X"82",X"64",X"72",X"95",X"AC",X"A3",X"A7",
		X"9E",X"90",X"77",X"69",X"82",X"AC",X"AC",X"8B",X"6E",X"43",X"56",X"72",X"99",X"B6",X"9E",X"80",
		X"5B",X"35",X"27",X"43",X"6E",X"90",X"95",X"77",X"4D",X"56",X"77",X"95",X"BF",X"D7",X"C8",X"9E",
		X"7C",X"5B",X"43",X"69",X"87",X"A7",X"B6",X"8B",X"72",X"4D",X"51",X"77",X"90",X"B6",X"A3",X"80",
		X"60",X"43",X"64",X"82",X"A3",X"C4",X"DB",X"CD",X"B1",X"8B",X"8B",X"AC",X"CD",X"D2",X"BA",X"99",
		X"77",X"5B",X"72",X"90",X"B6",X"C4",X"A7",X"82",X"7C",X"9E",X"BF",X"BA",X"95",X"9E",X"99",X"99",
		X"A3",X"9E",X"9E",X"99",X"95",X"99",X"9E",X"AC",X"B6",X"9E",X"87",X"64",X"64",X"82",X"A3",X"B1",
		X"9E",X"80",X"5B",X"43",X"5B",X"7C",X"9E",X"AC",X"90",X"6E",X"64",X"87",X"A7",X"B1",X"AC",X"99",
		X"7C",X"5B",X"3F",X"51",X"72",X"90",X"A7",X"8B",X"6E",X"48",X"43",X"60",X"82",X"87",X"60",X"43",
		X"1E",X"2C",X"56",X"77",X"90",X"77",X"5B",X"35",X"27",X"48",X"69",X"87",X"B1",X"AC",X"8B",X"69",
		X"43",X"56",X"72",X"69",X"6E",X"69",X"5B",X"4D",X"60",X"69",X"60",X"6E",X"80",X"82",X"6E",X"4D",
		X"56",X"5B",X"3F",X"27",X"35",X"60",X"72",X"69",X"6E",X"69",X"56",X"51",X"60",X"80",X"82",X"60",
		X"43",X"22",X"31",X"51",X"72",X"90",X"7C",X"60",X"3A",X"2C",X"35",X"31",X"3A",X"51",X"56",X"43",
		X"27",X"2C",X"51",X"6E",X"95",X"B6",X"9E",X"80",X"56",X"43",X"64",X"80",X"AC",X"B1",X"90",X"72",
		X"48",X"51",X"6E",X"90",X"B6",X"A3",X"82",X"60",X"43",X"60",X"7C",X"A7",X"B6",X"95",X"77",X"4D",
		X"4D",X"6E",X"90",X"8B",X"8B",X"8B",X"80",X"82",X"90",X"9E",X"95",X"77",X"69",X"80",X"AC",X"AC",
		X"A3",X"AC",X"99",X"8B",X"69",X"77",X"99",X"B6",X"A7",X"80",X"5B",X"48",X"60",X"82",X"AC",X"B6",
		X"95",X"6E",X"51",X"2C",X"31",X"5B",X"7C",X"99",X"8B",X"64",X"4D",X"60",X"87",X"A7",X"C8",X"DB",
		X"B6",X"90",X"77",X"51",X"51",X"77",X"90",X"B1",X"A7",X"82",X"64",X"48",X"64",X"80",X"A3",X"B6",
		X"95",X"77",X"4D",X"51",X"72",X"90",X"BA",X"D7",X"DB",X"C4",X"99",X"82",X"95",X"BF",X"D7",X"CD",
		X"B1",X"87",X"64",X"60",X"82",X"A7",X"C8",X"BF",X"99",X"77",X"87",X"A7",X"C4",X"A7",X"95",X"A3",
		X"99",X"A7",X"A3",X"A3",X"9E",X"99",X"99",X"9E",X"A7",X"BA",X"B1",X"99",X"72",X"60",X"72",X"99",
		X"B6",X"B1",X"95",X"6E",X"4D",X"48",X"6E",X"90",X"B1",X"A7",X"80",X"60",X"77",X"95",X"B1",X"B1",
		X"AC",X"95",X"6E",X"48",X"3F",X"64",X"87",X"A7",X"A3",X"82",X"5B",X"3F",X"4D",X"77",X"90",X"77",
		X"5B",X"31",X"22",X"43",X"60",X"8B",X"8B",X"6E",X"4D",X"27",X"35",X"56",X"77",X"9E",X"B6",X"A3",
		X"7C",X"5B",X"43",X"69",X"72",X"69",X"72",X"64",X"51",X"51",X"69",X"69",X"69",X"77",X"82",X"80",
		X"60",X"51",X"60",X"51",X"35",X"2C",X"48",X"77",X"72",X"6E",X"72",X"64",X"56",X"56",X"72",X"8B",
		X"7C",X"5B",X"35",X"1E",X"3F",X"5B",X"8B",X"90",X"72",X"51",X"27",X"35",X"35",X"35",X"48",X"56",
		X"56",X"35",X"22",X"3A",X"60",X"82",X"A7",X"B1",X"95",X"6E",X"4D",X"4D",X"72",X"95",X"B6",X"A3",
		X"80",X"60",X"43",X"64",X"82",X"A3",X"B6",X"90",X"77",X"51",X"4D",X"77",X"90",X"B6",X"A7",X"82",
		X"64",X"48",X"5B",X"82",X"95",X"87",X"8B",X"82",X"82",X"87",X"9E",X"9E",X"8B",X"72",X"72",X"95",
		X"B1",X"A7",X"A7",X"A3",X"99",X"7C",X"69",X"82",X"A3",X"B6",X"90",X"77",X"51",X"51",X"77",X"90",
		X"B1",X"A7",X"82",X"69",X"3F",X"27",X"48",X"64",X"90",X"99",X"7C",X"5B",X"56",X"77",X"90",X"B6",
		X"DB",X"CD",X"A7",X"87",X"60",X"48",X"60",X"82",X"A7",X"B6",X"99",X"77",X"51",X"4D",X"72",X"95",
		X"B6",X"AC",X"87",X"64",X"48",X"5B",X"82",X"A3",X"C4",X"DB",X"D2",X"B6",X"90",X"87",X"AC",X"CD",
		X"D7",X"C4",X"9E",X"80",X"60",X"72",X"95",X"B6",X"CD",X"AC",X"87",X"7C",X"95",X"BF",X"C4",X"99",
		X"99",X"9E",X"9E",X"A7",X"A3",X"A3",X"9E",X"99",X"99",X"A3",X"AC",X"BA",X"A7",X"8B",X"69",X"60",
		X"87",X"A3",X"B6",X"A7",X"82",X"64",X"43",X"5B",X"7C",X"9E",X"B6",X"95",X"72",X"64",X"80",X"A7",
		X"B6",X"B1",X"A7",X"80",X"64",X"3F",X"4D",X"77",X"90",X"B1",X"95",X"77",X"51",X"43",X"60",X"82",
		X"8B",X"64",X"48",X"22",X"2C",X"56",X"77",X"95",X"80",X"5B",X"3F",X"22",X"48",X"69",X"87",X"A7",
		X"B1",X"90",X"72",X"4D",X"51",X"77",X"6E",X"6E",X"6E",X"60",X"4D",X"60",X"6E",X"64",X"6E",X"80",
		X"82",X"77",X"5B",X"56",X"5B",X"48",X"31",X"35",X"60",X"77",X"6E",X"72",X"6E",X"60",X"56",X"60",
		X"80",X"8B",X"64",X"48",X"27",X"27",X"56",X"6E",X"95",X"80",X"60",X"3F",X"27",X"35",X"35",X"3A",
		X"4D",X"56",X"48",X"2C",X"27",X"51",X"72",X"90",X"B1",X"A3",X"82",X"64",X"48",X"60",X"80",X"9E",
		X"B1",X"95",X"77",X"51",X"4D",X"72",X"8B",X"B1",X"A7",X"87",X"69",X"48",X"5B",X"80",X"9E",X"B6",
		X"99",X"7C",X"56",X"4D",X"69",X"90",X"90",X"8B",X"8B",X"80",X"82",X"90",X"9E",X"99",X"7C",X"69",
		X"80",X"A3",X"AC",X"A3",X"AC",X"9E",X"90",X"6E",X"72",X"90",X"B6",X"A7",X"87",X"64",X"43",X"60",
		X"7C",X"A7",X"B6",X"99",X"7C",X"56",X"31",X"31",X"51",X"7C",X"99",X"90",X"6E",X"4D",X"60",X"80",
		X"A3",X"CD",X"DB",X"C4",X"95",X"7C",X"56",X"4D",X"77",X"90",X"B6",X"AC",X"87",X"69",X"48",X"48",
		X"48",X"43",X"48",X"51",X"5B",X"51",X"4D",X"5B",X"5B",X"51",X"56",X"60",X"60",X"51",X"43",X"4D",
		X"60",X"87",X"AC",X"BF",X"A3",X"7C",X"56",X"51",X"72",X"95",X"BA",X"B6",X"90",X"6E",X"7C",X"99",
		X"8B",X"95",X"A3",X"99",X"7C",X"6E",X"87",X"AC",X"B1",X"95",X"72",X"72",X"77",X"77",X"77",X"6E",
		X"77",X"7C",X"77",X"72",X"77",X"7C",X"8B",X"95",X"82",X"6E",X"48",X"48",X"69",X"87",X"A7",X"9E",
		X"80",X"60",X"43",X"56",X"77",X"99",X"AC",X"90",X"72",X"51",X"48",X"69",X"87",X"AC",X"A7",X"82",
		X"64",X"48",X"56",X"77",X"99",X"B1",X"99",X"77",X"5B",X"31",X"2C",X"4D",X"6E",X"95",X"90",X"72",
		X"51",X"5B",X"80",X"99",X"BA",X"A3",X"82",X"60",X"4D",X"6E",X"8B",X"AC",X"B6",X"90",X"77",X"51",
		X"5B",X"7C",X"99",X"8B",X"69",X"82",X"9E",X"80",X"6E",X"8B",X"A3",X"D2",X"D7",X"B6",X"90",X"90",
		X"B1",X"CD",X"EE",X"E0",X"BF",X"99",X"80",X"90",X"B6",X"CD",X"AC",X"87",X"6E",X"48",X"43",X"64",
		X"87",X"82",X"5B",X"6E",X"69",X"56",X"60",X"77",X"90",X"72",X"64",X"72",X"60",X"43",X"3F",X"64",
		X"87",X"82",X"60",X"43",X"4D",X"77",X"8B",X"BA",X"CD",X"B1",X"95",X"69",X"60",X"7C",X"9E",X"A3",
		X"82",X"64",X"43",X"1E",X"31",X"51",X"77",X"95",X"80",X"60",X"48",X"64",X"82",X"A7",X"AC",X"90",
		X"6E",X"6E",X"77",X"5B",X"64",X"77",X"72",X"60",X"69",X"80",X"A7",X"B6",X"9E",X"77",X"69",X"8B",
		X"90",X"87",X"9E",X"9E",X"8B",X"64",X"4D",X"56",X"80",X"99",X"87",X"90",X"87",X"7C",X"64",X"3F",
		X"3A",X"56",X"7C",X"80",X"56",X"3A",X"43",X"69",X"8B",X"AC",X"C8",X"AC",X"8B",X"69",X"56",X"7C",
		X"99",X"A3",X"80",X"80",X"99",X"BF",X"BA",X"90",X"A3",X"BF",X"AC",X"8B",X"A7",X"BF",X"A3",X"7C",
		X"6E",X"87",X"B1",X"CD",X"F3",X"F3",X"C4",X"A7",X"82",X"90",X"B6",X"D2",X"EE",X"D2",X"AC",X"95",
		X"B6",X"BF",X"B1",X"C8",X"C8",X"B1",X"95",X"95",X"BA",X"DB",X"C8",X"A3",X"8B",X"95",X"8B",X"90",
		X"8B",X"87",X"8B",X"90",X"87",X"87",X"8B",X"95",X"A7",X"A3",X"90",X"6E",X"4D",X"64",X"80",X"A7",
		X"BF",X"9E",X"82",X"56",X"4D",X"72",X"95",X"B6",X"B1",X"8B",X"64",X"48",X"5B",X"80",X"A3",X"BA",
		X"9E",X"7C",X"56",X"48",X"69",X"8B",X"B1",X"B1",X"8B",X"64",X"48",X"27",X"3A",X"60",X"80",X"99",
		X"80",X"5B",X"48",X"69",X"8B",X"B1",X"B6",X"90",X"6E",X"4D",X"51",X"77",X"99",X"B6",X"A3",X"80",
		X"5B",X"48",X"60",X"87",X"95",X"72",X"69",X"90",X"90",X"69",X"72",X"95",X"B1",X"C8",X"B6",X"8B",
		X"77",X"87",X"B1",X"C8",X"BF",X"A3",X"7C",X"5B",X"56",X"77",X"9E",X"95",X"77",X"51",X"2C",X"14",
		X"22",X"4D",X"69",X"4D",X"3A",X"48",X"35",X"31",X"43",X"69",X"69",X"43",X"4D",X"4D",X"3A",X"1E",
		X"2C",X"5B",X"6E",X"60",X"31",X"22",X"3F",X"64",X"87",X"AC",X"AC",X"8B",X"69",X"48",X"4D",X"77",
		X"95",X"82",X"64",X"3F",X"19",X"0B",X"27",X"4D",X"77",X"7C",X"60",X"35",X"3A",X"5B",X"80",X"A3",
		X"90",X"72",X"56",X"64",X"5B",X"48",X"60",X"69",X"56",X"4D",X"64",X"7C",X"A3",X"A3",X"7C",X"5B",
		X"64",X"82",X"7C",X"82",X"95",X"87",X"72",X"4D",X"3F",X"60",X"82",X"87",X"80",X"82",X"77",X"6E",
		X"48",X"27",X"35",X"64",X"7C",X"64",X"43",X"31",X"4D",X"72",X"8B",X"BA",X"BA",X"99",X"7C",X"51",
		X"60",X"7C",X"99",X"8B",X"72",X"82",X"A7",X"BF",X"9E",X"8B",X"B1",X"BA",X"95",X"8B",X"B6",X"B1",
		X"8B",X"6E",X"77",X"99",X"B6",X"DB",X"F7",X"D7",X"BA",X"8B",X"80",X"9E",X"BA",X"E5",X"E5",X"BF",
		X"9E",X"9E",X"C4",X"B1",X"BA",X"C8",X"BF",X"A3",X"8B",X"A3",X"C8",X"D7",X"B6",X"8B",X"87",X"90",
		X"8B",X"90",X"87",X"87",X"8B",X"8B",X"82",X"87",X"8B",X"99",X"A7",X"95",X"80",X"5B",X"4D",X"77",
		X"90",X"B6",X"B1",X"87",X"6E",X"48",X"5B",X"82",X"9E",X"BA",X"9E",X"7C",X"5B",X"48",X"6E",X"8B",
		X"B1",X"B1",X"87",X"6E",X"48",X"56",X"7C",X"99",X"B6",X"9E",X"7C",X"60",X"3A",X"2C",X"48",X"69",
		X"8B",X"90",X"72",X"51",X"51",X"7C",X"95",X"BA",X"A3",X"80",X"64",X"43",X"64",X"82",X"A7",X"B6",
		X"90",X"77",X"4D",X"4D",X"72",X"90",X"8B",X"69",X"7C",X"95",X"82",X"69",X"80",X"9E",X"BA",X"BF",
		X"A3",X"80",X"77",X"99",X"BA",X"C4",X"B1",X"8B",X"6E",X"4D",X"60",X"87",X"9E",X"82",X"5B",X"43",
		X"1E",X"14",X"35",X"5B",X"60",X"35",X"43",X"43",X"31",X"3A",X"4D",X"72",X"51",X"3F",X"51",X"48",
		X"22",X"1E",X"3F",X"60",X"69",X"48",X"27",X"2C",X"56",X"72",X"95",X"B1",X"9E",X"7C",X"5B",X"48",
		X"60",X"82",X"90",X"72",X"51",X"31",X"10",X"14",X"3A",X"5B",X"7C",X"6E",X"4D",X"31",X"4D",X"6E",
		X"90",X"A3",X"82",X"60",X"5B",X"69",X"4D",X"51",X"64",X"64",X"4D",X"5B",X"69",X"90",X"AC",X"90",
		X"72",X"5B",X"80",X"87",X"7C",X"90",X"90",X"82",X"64",X"3F",X"48",X"6E",X"87",X"80",X"82",X"82",
		X"72",X"60",X"3A",X"27",X"4D",X"72",X"7C",X"5B",X"31",X"3A",X"5B",X"80",X"A3",X"BF",X"B1",X"8B",
		X"64",X"51",X"69",X"90",X"A3",X"80",X"77",X"95",X"BA",X"BA",X"95",X"99",X"BA",X"B1",X"8B",X"9E",
		X"BA",X"A7",X"7C",X"69",X"82",X"A3",X"C8",X"EE",X"F3",X"CD",X"A7",X"82",X"87",X"A7",X"D2",X"E9",
		X"DB",X"B1",X"90",X"B1",X"C4",X"B1",X"C4",X"C8",X"BA",X"95",X"90",X"B1",X"D2",X"CD",X"A7",X"87",
		X"90",X"90",X"90",X"8B",X"87",X"8B",X"90",X"8B",X"87",X"8B",X"90",X"A7",X"A3",X"90",X"72",X"4D",
		X"64",X"80",X"A7",X"BF",X"A3",X"82",X"5B",X"4D",X"6E",X"87",X"B6",X"B1",X"90",X"72",X"48",X"5B",
		X"77",X"99",X"BA",X"9E",X"82",X"5B",X"48",X"69",X"82",X"B1",X"B1",X"90",X"72",X"48",X"2C",X"31",
		X"56",X"80",X"99",X"87",X"60",X"48",X"64",X"80",X"AC",X"B6",X"95",X"7C",X"4D",X"51",X"72",X"90",
		X"BA",X"A7",X"87",X"64",X"43",X"60",X"80",X"95",X"77",X"69",X"87",X"90",X"6E",X"6E",X"8B",X"B1",
		X"C8",X"BA",X"95",X"72",X"87",X"A3",X"C4",X"BF",X"A3",X"87",X"5B",X"51",X"72",X"90",X"95",X"77",
		X"5B",X"35",X"10",X"22",X"43",X"64",X"51",X"35",X"4D",X"3A",X"31",X"43",X"60",X"6E",X"48",X"48",
		X"51",X"3A",X"1E",X"22",X"51",X"72",X"60",X"3A",X"27",X"3F",X"64",X"80",X"AC",X"B1",X"90",X"72",
		X"48",X"4D",X"6E",X"90",X"87",X"64",X"48",X"22",X"06",X"27",X"43",X"72",X"80",X"64",X"43",X"3A",
		X"5B",X"7C",X"9E",X"99",X"77",X"56",X"64",X"60",X"4D",X"5B",X"69",X"60",X"51",X"60",X"7C",X"A3",
		X"A7",X"87",X"60",X"64",X"87",X"82",X"82",X"99",X"8B",X"77",X"51",X"3F",X"5B",X"82",X"8B",X"80",
		X"87",X"7C",X"72",X"51",X"2C",X"35",X"5B",X"7C",X"6E",X"48",X"31",X"4D",X"72",X"8B",X"B1",X"BA",
		X"9E",X"80",X"5B",X"5B",X"7C",X"9E",X"95",X"95",X"AC",X"C8",X"E5",X"CD",X"AC",X"87",X"77",X"90",
		X"B1",X"D7",X"D7",X"B6",X"90",X"95",X"BA",X"D7",X"C8",X"A7",X"B6",X"AC",X"B1",X"B6",X"B1",X"B1",
		X"AC",X"A7",X"AC",X"B1",X"C4",X"C4",X"AC",X"90",X"72",X"7C",X"99",X"BA",X"D7",X"BF",X"99",X"7C",
		X"69",X"82",X"A3",X"C8",X"C8",X"A7",X"82",X"87",X"AC",X"C8",X"D2",X"CD",X"B6",X"90",X"72",X"5B",
		X"77",X"90",X"B6",X"BF",X"9E",X"82",X"60",X"60",X"80",X"9E",X"95",X"6E",X"51",X"31",X"4D",X"72",
		X"90",X"A7",X"82",X"64",X"43",X"3A",X"60",X"80",X"9E",X"BF",X"B6",X"90",X"77",X"56",X"6E",X"82",
		X"77",X"7C",X"72",X"64",X"5B",X"72",X"72",X"6E",X"7C",X"8B",X"8B",X"77",X"5B",X"64",X"60",X"48",
		X"31",X"43",X"6E",X"7C",X"72",X"77",X"6E",X"60",X"5B",X"6E",X"8B",X"87",X"60",X"43",X"22",X"3A",
		X"60",X"80",X"99",X"7C",X"5B",X"35",X"31",X"3A",X"35",X"43",X"56",X"56",X"43",X"27",X"35",X"5B",
		X"77",X"A3",X"B6",X"99",X"7C",X"51",X"48",X"69",X"87",X"B1",X"AC",X"8B",X"69",X"43",X"56",X"77",
		X"99",X"B6",X"99",X"80",X"56",X"48",X"69",X"82",X"B1",X"AC",X"90",X"6E",X"48",X"51",X"77",X"90",
		X"87",X"8B",X"87",X"80",X"82",X"95",X"9E",X"8B",X"72",X"69",X"87",X"B1",X"A7",X"A3",X"A7",X"95",
		X"87",X"64",X"7C",X"9E",X"B6",X"9E",X"77",X"51",X"48",X"64",X"8B",X"AC",X"AC",X"8B",X"64",X"48",
		X"27",X"35",X"60",X"80",X"99",X"80",X"5B",X"4D",X"64",X"8B",X"AC",X"CD",X"D2",X"A7",X"8B",X"69",
		X"4D",X"56",X"77",X"95",X"B1",X"99",X"7C",X"5B",X"48",X"69",X"82",X"A7",X"AC",X"8B",X"6E",X"4D",
		X"51",X"77",X"90",X"B6",X"D7",X"D2",X"BF",X"90",X"80",X"99",X"BA",X"D2",X"C4",X"A7",X"87",X"5B",
		X"64",X"82",X"A7",X"C8",X"B6",X"90",X"77",X"8B",X"AC",X"C4",X"9E",X"95",X"9E",X"95",X"A3",X"9E",
		X"9E",X"9E",X"95",X"95",X"99",X"A7",X"B6",X"A7",X"95",X"6E",X"5B",X"77",X"95",X"B1",X"A7",X"8B",
		X"6E",X"43",X"4D",X"6E",X"95",X"AC",X"9E",X"77",X"60",X"77",X"99",X"B1",X"AC",X"A7",X"87",X"64",
		X"3F",X"43",X"69",X"8B",X"A7",X"99",X"77",X"51",X"3A",X"4D",X"7C",X"8B",X"6E",X"51",X"22",X"22",
		X"43",X"64",X"90",X"82",X"69",X"43",X"22",X"3A",X"56",X"80",X"A3",X"B6",X"99",X"72",X"51",X"43",
		X"6E",X"6E",X"69",X"6E",X"60",X"4D",X"56",X"69",X"64",X"69",X"77",X"82",X"77",X"5B",X"4D",X"60",
		X"48",X"2C",X"27",X"4D",X"77",X"6E",X"6E",X"6E",X"60",X"51",X"56",X"77",X"8B",X"72",X"56",X"27",
		X"22",X"43",X"64",X"90",X"87",X"6E",X"48",X"22",X"35",X"31",X"35",X"48",X"56",X"51",X"2C",X"22",
		X"3F",X"64",X"87",X"AC",X"AC",X"87",X"64",X"43",X"51",X"77",X"99",X"B1",X"9E",X"7C",X"56",X"43",
		X"60",X"87",X"AC",X"B1",X"90",X"69",X"48",X"4D",X"72",X"95",X"B6",X"A3",X"80",X"5B",X"48",X"5B",
		X"87",X"90",X"82",X"90",X"80",X"82",X"87",X"99",X"99",X"82",X"69",X"72",X"9E",X"B1",X"A3",X"A7",
		X"9E",X"95",X"7C",X"6E",X"87",X"AC",X"B1",X"87",X"6E",X"48",X"56",X"7C",X"95",X"B6",X"9E",X"7C",
		X"60",X"35",X"27",X"4D",X"69",X"95",X"95",X"77",X"56",X"56",X"7C",X"95",X"BF",X"DB",X"C4",X"A3",
		X"80",X"56",X"48",X"64",X"8B",X"AC",X"B1",X"90",X"6E",X"4D",X"51",X"77",X"99",X"B6",X"A7",X"80",
		X"5B",X"48",X"60",X"87",X"A7",X"C8",X"DB",X"CD",X"B1",X"87",X"8B",X"B1",X"CD",X"D7",X"BA",X"95",
		X"77",X"5B",X"7C",X"99",X"BA",X"C8",X"A3",X"82",X"7C",X"99",X"C4",X"BA",X"95",X"9E",X"99",X"9E",
		X"A7",X"A3",X"A3",X"9E",X"95",X"9E",X"A3",X"B1",X"BA",X"9E",X"87",X"60",X"69",X"8B",X"A7",X"B6",
		X"9E",X"7C",X"5B",X"43",X"60",X"80",X"A3",X"B1",X"8B",X"6E",X"69",X"87",X"AC",X"B1",X"B1",X"9E",
		X"77",X"5B",X"3A",X"56",X"7C",X"99",X"B1",X"8B",X"6E",X"48",X"43",X"69",X"87",X"87",X"64",X"3F",
		X"22",X"31",X"56",X"80",X"95",X"80",X"5B",X"31",X"27",X"43",X"6E",X"8B",X"B1",X"B1",X"87",X"6E",
		X"43",X"56",X"77",X"69",X"72",X"69",X"5B",X"4D",X"60",X"69",X"64",X"6E",X"80",X"82",X"72",X"51",
		X"56",X"5B",X"43",X"27",X"3A",X"69",X"77",X"6E",X"6E",X"6E",X"5B",X"51",X"64",X"82",X"87",X"60",
		X"43",X"1E",X"31",X"5B",X"77",X"95",X"7C",X"5B",X"35",X"2C",X"35",X"35",X"3F",X"51",X"56",X"43",
		X"27",X"2C",X"5B",X"77",X"95",X"B1",X"9E",X"7C",X"5B",X"48",X"69",X"82",X"A7",X"AC",X"8B",X"72",
		X"4D",X"51",X"77",X"95",X"B1",X"A3",X"80",X"60",X"48",X"64",X"82",X"A3",X"B1",X"90",X"77",X"51",
		X"51",X"72",X"95",X"8B",X"8B",X"8B",X"80",X"87",X"95",X"9E",X"95",X"77",X"69",X"82",X"A7",X"AC",
		X"A7",X"AC",X"99",X"87",X"6E",X"77",X"99",X"BA",X"9E",X"82",X"5B",X"48",X"69",X"82",X"B1",X"B1",
		X"95",X"72",X"4D",X"2C",X"35",X"5B",X"80",X"99",X"8B",X"64",X"4D",X"69",X"87",X"AC",X"D2",X"D7",
		X"BA",X"90",X"72",X"4D",X"51",X"7C",X"95",X"BA",X"A7",X"82",X"64",X"48",X"69",X"87",X"A7",X"BA",
		X"90",X"77",X"51",X"51",X"77",X"95",X"B1",X"D7",X"DB",X"C4",X"A3",X"87",X"99",X"BF",X"D7",X"CD",
		X"AC",X"8B",X"69",X"64",X"87",X"A3",X"C8",X"BA",X"99",X"7C",X"8B",X"B1",X"C8",X"AC",X"99",X"A3",
		X"99",X"A3",X"A3",X"A3",X"A3",X"99",X"99",X"9E",X"A3",X"B6",X"AC",X"99",X"72",X"5B",X"77",X"95",
		X"B6",X"B1",X"90",X"72",X"48",X"4D",X"6E",X"8B",X"B6",X"A3",X"82",X"64",X"77",X"99",X"B1",X"B1",
		X"A7",X"90",X"72",X"43",X"43",X"64",X"82",X"AC",X"9E",X"82",X"5B",X"3A",X"51",X"72",X"8B",X"77",
		X"56",X"35",X"22",X"48",X"64",X"87",X"8B",X"6E",X"4D",X"2C",X"35",X"5B",X"77",X"9E",X"BA",X"9E",
		X"80",X"56",X"43",X"6E",X"72",X"6E",X"6E",X"64",X"56",X"56",X"6E",X"64",X"69",X"77",X"82",X"80",
		X"60",X"51",X"60",X"51",X"31",X"2C",X"4D",X"6E",X"72",X"6E",X"72",X"64",X"51",X"5B",X"72",X"87",
		X"77",X"56",X"35",X"22",X"43",X"60",X"87",X"8B",X"6E",X"51",X"2C",X"35",X"35",X"35",X"48",X"56",
		X"51",X"3A",X"27",X"3F",X"64",X"80",X"AC",X"B1",X"90",X"72",X"48",X"51",X"72",X"90",X"B6",X"A3",
		X"87",X"60",X"43",X"60",X"80",X"A7",X"B6",X"95",X"77",X"4D",X"4D",X"72",X"90",X"BA",X"A7",X"8B",
		X"64",X"48",X"5B",X"80",X"95",X"87",X"90",X"82",X"82",X"87",X"99",X"9E",X"87",X"6E",X"6E",X"95",
		X"B6",X"A3",X"AC",X"A3",X"95",X"80",X"69",X"87",X"AC",X"B6",X"8B",X"72",X"4D",X"51",X"7C",X"95",
		X"BA",X"A3",X"80",X"64",X"43",X"2C",X"48",X"69",X"8B",X"95",X"7C",X"56",X"51",X"7C",X"95",X"BA",
		X"D7",X"C8",X"A3",X"87",X"60",X"48",X"64",X"80",X"AC",X"B6",X"95",X"77",X"4D",X"48",X"48",X"48",
		X"4D",X"4D",X"4D",X"51",X"51",X"51",X"51",X"56",X"56",X"56",X"56",X"5B",X"5B",X"5B",X"5B",X"5B",
		X"60",X"60",X"60",X"60",X"60",X"64",X"64",X"64",X"64",X"64",X"64",X"69",X"69",X"69",X"69",X"69",
		X"69",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"6E",X"72",X"72",X"72",X"72",X"72",X"72",X"72",X"72",
		X"72",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"77",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"82",X"82",X"87",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",
		X"80",X"80",X"80",X"80",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"80",X"7C",X"7C",
		X"7C",X"7C",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"7C",
		X"80",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"7C",
		X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"80",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"80",X"80",X"7C",X"77",X"77",X"7C",X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"7C",X"80",X"82",
		X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"77",X"7C",
		X"7C",X"80",X"82",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",
		X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",
		X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"82",X"7C",X"7C",
		X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",
		X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"72",X"77",X"80",X"82",X"7C",X"77",X"82",X"82",X"7C",X"7C",
		X"82",X"82",X"77",X"7C",X"82",X"80",X"77",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",
		X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",
		X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",
		X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",
		X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",
		X"7C",X"77",X"72",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",
		X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"82",X"80",X"7C",X"7C",X"82",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"72",X"77",X"7C",X"7C",X"7C",X"7C",X"80",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",
		X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"82",X"80",
		X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",
		X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",
		X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",
		X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"80",X"80",X"77",X"7C",X"80",X"7C",X"77",X"7C",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"82",X"82",X"77",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",
		X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",
		X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"72",X"77",X"7C",X"7C",X"7C",X"7C",X"77",X"7C",X"7C",X"7C",X"7C",
		X"77",X"77",X"7C",X"7C",X"77",X"77",X"7C",X"7C",X"80",X"7C",X"7C",X"7C",X"80",X"7C",X"82",X"82",
		X"80",X"7C",X"7C",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",
		X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"82",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"82",X"82",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"80",
		X"7C",X"80",X"87",X"87",X"87",X"8B",X"8B",X"8B",X"95",X"90",X"90",X"99",X"95",X"95",X"95",X"95",
		X"90",X"95",X"99",X"95",X"87",X"87",X"8B",X"82",X"7C",X"7C",X"80",X"77",X"6E",X"72",X"72",X"69",
		X"64",X"69",X"60",X"5B",X"48",X"48",X"4D",X"48",X"56",X"51",X"4D",X"51",X"51",X"51",X"5B",X"64",
		X"60",X"64",X"69",X"69",X"72",X"72",X"72",X"77",X"80",X"80",X"80",X"87",X"8B",X"87",X"8B",X"95",
		X"99",X"90",X"99",X"99",X"95",X"90",X"95",X"95",X"90",X"87",X"87",X"87",X"80",X"7C",X"80",X"7C",
		X"77",X"77",X"72",X"72",X"72",X"6E",X"69",X"72",X"7C",X"7C",X"6E",X"72",X"7C",X"7C",X"7C",X"82",
		X"87",X"82",X"7C",X"82",X"87",X"82",X"87",X"8B",X"82",X"82",X"82",X"80",X"80",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"80",X"7C",X"82",X"82",X"82",X"82",X"82",X"87",X"87",X"87",X"87",X"87",
		X"87",X"80",X"82",X"87",X"82",X"87",X"8B",X"87",X"80",X"7C",X"87",X"87",X"7C",X"80",X"80",X"77",
		X"7C",X"7C",X"7C",X"77",X"7C",X"80",X"7C",X"7C",X"7C",X"72",X"72",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"72",X"77",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"72",X"7C",X"7C",X"7C",X"82",
		X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",
		X"80",X"80",X"82",X"80",X"77",X"80",X"82",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"77",X"72",X"77",X"7C",X"77",X"72",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"72",X"77",X"7C",X"7C",X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"80",X"77",X"77",
		X"77",X"77",X"77",X"77",X"80",X"87",X"80",X"77",X"80",X"7C",X"77",X"7C",X"82",X"82",X"82",X"82",
		X"80",X"77",X"77",X"80",X"90",X"87",X"77",X"80",X"7C",X"80",X"82",X"80",X"87",X"87",X"82",X"7C",
		X"77",X"82",X"80",X"80",X"87",X"82",X"80",X"77",X"7C",X"7C",X"80",X"82",X"80",X"82",X"7C",X"7C",
		X"7C",X"77",X"72",X"7C",X"82",X"80",X"77",X"7C",X"7C",X"72",X"77",X"80",X"82",X"7C",X"77",X"7C",
		X"77",X"77",X"7C",X"82",X"82",X"77",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"82",X"7C",X"7C",
		X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"77",X"77",X"7C",X"7C",X"80",X"7C",X"77",X"77",X"77",X"7C",X"80",X"7C",
		X"7C",X"7C",X"80",X"77",X"77",X"80",X"80",X"80",X"7C",X"77",X"7C",X"80",X"87",X"80",X"7C",X"82",
		X"87",X"80",X"7C",X"82",X"82",X"82",X"82",X"82",X"82",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",
		X"80",X"82",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"82",X"80",X"7C",X"7C",X"82",X"80",
		X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"77",X"6E",X"77",X"80",X"7C",
		X"80",X"82",X"80",X"72",X"72",X"7C",X"80",X"72",X"72",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"72",
		X"7C",X"80",X"77",X"72",X"7C",X"7C",X"7C",X"82",X"82",X"7C",X"72",X"77",X"80",X"7C",X"80",X"82",
		X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"82",X"80",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"80",X"82",X"80",X"82",X"80",X"7C",X"82",X"82",X"80",X"80",X"7C",X"7C",X"7C",
		X"80",X"82",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"82",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"82",X"7C",X"7C",X"7C",X"7C",X"82",
		X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"77",X"72",X"80",X"7C",X"7C",
		X"82",X"80",X"7C",X"72",X"7C",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",
		X"80",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"82",X"80",
		X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",
		X"80",X"7C",X"7C",X"7C",X"72",X"77",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"77",X"77",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",
		X"80",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",
		X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",
		X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",
		X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"7C",X"7C",X"80",X"82",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"82",X"80",X"7C",X"80",
		X"80",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",
		X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"80",X"82",
		X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",
		X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"77",X"7C",X"82",
		X"7C",X"77",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",
		X"77",X"7C",X"82",X"7C",X"77",X"80",X"80",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"80",X"80",X"77",
		X"7C",X"82",X"7C",X"77",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"82",X"7C",X"7C",
		X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",
		X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",
		X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",
		X"80",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",
		X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"80",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",
		X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",X"7C",X"80",
		X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",
		X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",
		X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",X"80",
		X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"82",X"80",X"7C",X"80",X"82",
		X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"77",X"7C",X"82",X"7C",
		X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",
		X"82",X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"82",X"80",X"7C",X"7C",X"82",
		X"80",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",
		X"7C",X"80",X"82",X"7C",X"7C",X"80",X"82",X"7C",X"7C",X"80",X"80",X"7C",X"7C",X"82",X"80",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"80",X"82",X"80",X"7C",X"80",
		X"82",X"8B",X"82",X"7C",X"87",X"87",X"80",X"80",X"87",X"87",X"80",X"6E",X"6E",X"87",X"A3",X"C4",
		X"E0",X"C8",X"A3",X"82",X"6E",X"8B",X"A7",X"CD",X"D2",X"B1",X"8B",X"8B",X"B6",X"A3",X"A7",X"B6",
		X"B1",X"95",X"80",X"95",X"BA",X"C8",X"B1",X"80",X"80",X"87",X"80",X"82",X"7C",X"80",X"82",X"82",
		X"7C",X"80",X"82",X"90",X"9E",X"90",X"77",X"51",X"43",X"64",X"87",X"AC",X"AC",X"87",X"64",X"43",
		X"4D",X"77",X"99",X"B1",X"9E",X"77",X"51",X"43",X"60",X"82",X"A7",X"AC",X"8B",X"64",X"43",X"4D",
		X"6E",X"95",X"B1",X"9E",X"7C",X"56",X"35",X"1E",X"43",X"64",X"87",X"8B",X"6E",X"4D",X"4D",X"77",
		X"90",X"B6",X"A3",X"7C",X"60",X"43",X"60",X"80",X"A3",X"B6",X"8B",X"72",X"4D",X"48",X"72",X"90",
		X"8B",X"69",X"77",X"90",X"80",X"64",X"7C",X"99",X"BF",X"CD",X"AC",X"87",X"80",X"A3",X"BF",X"E5",
		X"DB",X"B1",X"90",X"72",X"80",X"A7",X"BA",X"A7",X"80",X"60",X"3A",X"2C",X"51",X"77",X"7C",X"5B",
		X"5B",X"60",X"48",X"51",X"64",X"82",X"6E",X"5B",X"64",X"5B",X"3F",X"31",X"4D",X"72",X"7C",X"56",
		X"35",X"3A",X"5B",X"82",X"9E",X"C4",X"AC",X"87",X"69",X"4D",X"6E",X"90",X"9E",X"82",X"5B",X"3A",
		X"19",X"19",X"43",X"60",X"82",X"7C",X"51",X"3A",X"4D",X"72",X"95",X"A7",X"90",X"64",X"60",X"6E",
		X"56",X"56",X"69",X"6E",X"56",X"5B",X"6E",X"8B",X"AC",X"95",X"77",X"5B",X"80",X"8B",X"7C",X"8B",
		X"90",X"82",X"69",X"43",X"48",X"6E",X"8B",X"82",X"82",X"80",X"77",X"60",X"35",X"27",X"3F",X"72",
		X"77",X"5B",X"3A",X"35",X"5B",X"77",X"99",X"BF",X"AC",X"8B",X"69",X"4D",X"64",X"87",X"99",X"7C",
		X"72",X"8B",X"B6",X"B6",X"90",X"90",X"B6",X"AC",X"87",X"99",X"B6",X"A3",X"77",X"64",X"80",X"9E",
		X"C4",X"E5",X"EE",X"C8",X"9E",X"80",X"82",X"A3",X"C8",X"E5",X"D7",X"A7",X"8B",X"A7",X"BA",X"AC",
		X"BF",X"C4",X"B1",X"8B",X"8B",X"AC",X"CD",X"C8",X"9E",X"82",X"87",X"87",X"87",X"87",X"80",X"87",
		X"87",X"82",X"80",X"87",X"8B",X"9E",X"9E",X"8B",X"6E",X"4D",X"5B",X"7C",X"99",X"B6",X"9E",X"80",
		X"5B",X"48",X"69",X"82",X"A7",X"AC",X"8B",X"6E",X"4D",X"51",X"72",X"90",X"B1",X"9E",X"7C",X"5B",
		X"43",X"60",X"80",X"A3",X"AC",X"8B",X"6E",X"4D",X"22",X"2C",X"4D",X"72",X"95",X"82",X"64",X"48",
		X"60",X"80",X"9E",X"B1",X"90",X"72",X"51",X"4D",X"6E",X"87",X"AC",X"A3",X"82",X"64",X"43",X"56",
		X"7C",X"95",X"77",X"64",X"82",X"90",X"69",X"69",X"82",X"A3",X"C4",X"B6",X"95",X"77",X"80",X"A3",
		X"BF",X"BA",X"9E",X"82",X"5B",X"51",X"69",X"8B",X"95",X"72",X"51",X"35",X"10",X"1E",X"3F",X"64",
		X"4D",X"31",X"48",X"3A",X"31",X"3A",X"5B",X"6E",X"43",X"43",X"4D",X"3A",X"19",X"22",X"48",X"64",
		X"5B",X"35",X"1E",X"35",X"60",X"7C",X"A7",X"AC",X"8B",X"6E",X"43",X"48",X"6E",X"8B",X"82",X"60",
		X"48",X"1E",X"01",X"22",X"3F",X"6E",X"7C",X"60",X"3F",X"35",X"56",X"77",X"99",X"95",X"77",X"56",
		X"60",X"5B",X"48",X"56",X"64",X"5B",X"4D",X"5B",X"77",X"9E",X"A3",X"82",X"5B",X"60",X"82",X"80",
		X"80",X"95",X"87",X"77",X"4D",X"3A",X"51",X"80",X"87",X"7C",X"82",X"77",X"6E",X"51",X"2C",X"31",
		X"56",X"77",X"6E",X"43",X"2C",X"3F",X"69",X"8B",X"AC",X"BF",X"99",X"7C",X"56",X"51",X"7C",X"99",
		X"95",X"72",X"80",X"9E",X"BF",X"A7",X"87",X"A3",X"BA",X"99",X"87",X"AC",X"B6",X"90",X"6E",X"6E",
		X"8B",X"B6",X"D2",X"F3",X"E0",X"B6",X"99",X"7C",X"95",X"B6",X"DB",X"E9",X"C4",X"9E",X"95",X"BA",
		X"B6",X"B1",X"C8",X"C4",X"A7",X"8B",X"95",X"C4",X"D7",X"BF",X"99",X"87",X"90",X"8B",X"90",X"87",
		X"87",X"8B",X"8B",X"82",X"87",X"8B",X"95",X"A7",X"99",X"87",X"60",X"4D",X"6E",X"87",X"B6",X"B6",
		X"95",X"77",X"4D",X"56",X"77",X"95",X"BA",X"A3",X"87",X"60",X"48",X"64",X"80",X"AC",X"B6",X"95",
		X"72",X"4D",X"4D",X"72",X"99",X"B6",X"A7",X"82",X"60",X"3F",X"22",X"43",X"69",X"87",X"99",X"77",
		X"51",X"4D",X"72",X"95",X"B6",X"AC",X"87",X"64",X"48",X"5B",X"80",X"A3",X"B6",X"9E",X"77",X"51",
		X"48",X"69",X"90",X"90",X"69",X"72",X"95",X"87",X"69",X"7C",X"9E",X"BA",X"C8",X"A7",X"82",X"77",
		X"90",X"BA",X"C8",X"B6",X"99",X"72",X"51",X"56",X"80",X"9E",X"8B",X"6E",X"48",X"1E",X"10",X"2C",
		X"56",X"64",X"3F",X"3F",X"48",X"31",X"35",X"48",X"6E",X"60",X"3F",X"4D",X"48",X"31",X"19",X"35",
		X"60",X"6E",X"56",X"27",X"27",X"48",X"6E",X"90",X"B1",X"A7",X"82",X"5B",X"43",X"56",X"80",X"95",
		X"7C",X"5B",X"35",X"14",X"0B",X"31",X"56",X"7C",X"77",X"56",X"31",X"43",X"64",X"8B",X"A3",X"8B",
		X"6E",X"5B",X"69",X"56",X"4D",X"64",X"69",X"56",X"56",X"6E",X"87",X"AC",X"99",X"77",X"5B",X"72",
		X"87",X"7C",X"8B",X"95",X"82",X"6E",X"48",X"43",X"69",X"8B",X"82",X"80",X"82",X"77",X"69",X"3F",
		X"27",X"43",X"69",X"7C",X"60",X"3A",X"31",X"5B",X"7C",X"95",X"BA",X"B1",X"95",X"6E",X"51",X"69",
		X"87",X"9E",X"82",X"72",X"8B",X"B6",X"BF",X"95",X"95",X"BA",X"B6",X"8B",X"99",X"BA",X"A7",X"87",
		X"6E",X"80",X"A3",X"BF",X"E9",X"F3",X"D2",X"B1",X"82",X"87",X"A3",X"C4",X"EE",X"DB",X"BA",X"99",
		X"AC",X"C4",X"B1",X"C4",X"C8",X"BA",X"9E",X"90",X"AC",X"D2",X"D2",X"AC",X"87",X"90",X"90",X"90",
		X"90",X"87",X"8B",X"90",X"8B",X"82",X"8B",X"90",X"A3",X"A7",X"90",X"7C",X"51",X"5B",X"80",X"99",
		X"BF",X"A7",X"82",X"64",X"48",X"69",X"87",X"AC",X"BA",X"95",X"77",X"51",X"51",X"7C",X"95",X"B6",
		X"AC",X"82",X"69",X"48",X"64",X"82",X"A3",X"B6",X"95",X"77",X"56",X"35",X"31",X"51",X"72",X"95",
		X"8B",X"6E",X"4D",X"60",X"82",X"9E",X"BA",X"99",X"7C",X"5B",X"48",X"72",X"8B",X"B1",X"B1",X"87",
		X"6E",X"48",X"56",X"80",X"95",X"82",X"69",X"82",X"95",X"7C",X"6E",X"87",X"A7",X"C4",X"BA",X"9E",
		X"7C",X"80",X"A7",X"BF",X"C4",X"A7",X"87",X"64",X"4D",X"69",X"90",X"99",X"80",X"56",X"3A",X"14",
		X"19",X"43",X"64",X"5B",X"3A",X"48",X"3F",X"31",X"3F",X"5B",X"72",X"48",X"48",X"51",X"3F",X"1E",
		X"22",X"48",X"69",X"64",X"3F",X"22",X"35",X"60",X"7C",X"9E",X"B1",X"95",X"77",X"51",X"4D",X"6E",
		X"90",X"8B",X"69",X"4D",X"2C",X"0B",X"1E",X"43",X"64",X"80",X"69",X"43",X"31",X"5B",X"77",X"99",
		X"9E",X"7C",X"5B",X"60",X"64",X"4D",X"56",X"69",X"60",X"4D",X"60",X"72",X"9E",X"A7",X"8B",X"6E",
		X"60",X"87",X"82",X"80",X"99",X"8B",X"80",X"5B",X"3F",X"51",X"77",X"8B",X"80",X"87",X"80",X"72",
		X"56",X"31",X"31",X"5B",X"7C",X"77",X"51",X"31",X"43",X"64",X"87",X"B1",X"C4",X"A7",X"82",X"60",
		X"56",X"72",X"9E",X"99",X"90",X"A7",X"C8",X"E9",X"DB",X"B1",X"8B",X"72",X"87",X"AC",X"D2",X"E0",
		X"C4",X"95",X"90",X"B1",X"CD",X"D2",X"A7",X"B1",X"B1",X"B1",X"BA",X"B1",X"B6",X"AC",X"A7",X"AC",
		X"B1",X"C4",X"C8",X"B6",X"95",X"72",X"72",X"95",X"BA",X"D7",X"C8",X"A3",X"7C",X"64",X"7C",X"9E",
		X"C4",X"D2",X"B6",X"87",X"82",X"A3",X"C4",X"D2",X"CD",X"BF",X"99",X"77",X"5B",X"69",X"90",X"B6",
		X"C8",X"AC",X"82",X"60",X"56",X"77",X"9E",X"9E",X"7C",X"56",X"35",X"43",X"69",X"90",X"A7",X"90",
		X"69",X"43",X"3A",X"56",X"80",X"99",X"BF",X"BF",X"95",X"7C",X"51",X"64",X"82",X"72",X"7C",X"77",
		X"69",X"5B",X"6E",X"72",X"72",X"77",X"87",X"8B",X"7C",X"5B",X"60",X"64",X"48",X"31",X"3F",X"6E",
		X"80",X"72",X"77",X"72",X"60",X"5B",X"6E",X"87",X"8B",X"6E",X"48",X"27",X"31",X"56",X"80",X"99",
		X"82",X"60",X"3A",X"2C",X"3A",X"35",X"43",X"51",X"5B",X"48",X"27",X"2C",X"51",X"7C",X"95",X"B6",
		X"9E",X"7C",X"60",X"43",X"69",X"82",X"A7",X"B6",X"8B",X"72",X"4D",X"4D",X"77",X"90",X"B6",X"A3",
		X"80",X"64",X"43",X"64",X"82",X"A3",X"B6",X"90",X"77",X"4D",X"4D",X"72",X"95",X"8B",X"87",X"87",
		X"80",X"82",X"90",X"9E",X"95",X"7C",X"69",X"82",X"A7",X"AC",X"A3",X"A7",X"99",X"8B",X"69",X"77",
		X"95",X"B1",X"9E",X"80",X"60",X"48",X"64",X"80",X"A3",X"B1",X"90",X"72",X"51",X"27",X"31",X"51",
		X"77",X"99",X"87",X"69",X"4D",X"64",X"82",X"9E",X"CD",X"D7",X"B6",X"95",X"6E",X"4D",X"4D",X"72",
		X"95",X"B1",X"A7",X"82",X"60",X"43",X"60",X"82",X"A3",X"B6",X"8B",X"72",X"4D",X"4D",X"72",X"90",
		X"B1",X"D2",X"D7",X"BF",X"9E",X"82",X"95",X"BA",X"D2",X"C8",X"A7",X"8B",X"69",X"60",X"82",X"9E",
		X"C4",X"BA",X"95",X"77",X"87",X"AC",X"C4",X"A7",X"95",X"9E",X"95",X"A3",X"9E",X"9E",X"9E",X"95",
		X"95",X"99",X"A3",X"B6",X"AC",X"95",X"77",X"5B",X"72",X"95",X"AC",X"AC",X"8B",X"72",X"4D",X"48",
		X"6E",X"87",X"AC",X"A3",X"80",X"60",X"72",X"99",X"AC",X"B1",X"A7",X"8B",X"6E",X"4D",X"3F",X"64",
		X"80",X"A3",X"9E",X"80",X"60",X"3F",X"4D",X"72",X"8B",X"77",X"51",X"31",X"1E",X"43",X"60",X"87",
		X"8B",X"69",X"4D",X"27",X"31",X"56",X"77",X"95",X"B1",X"9E",X"7C",X"60",X"43",X"69",X"72",X"69",
		X"6E",X"64",X"51",X"51",X"69",X"64",X"64",X"77",X"82",X"7C",X"64",X"51",X"5B",X"51",X"35",X"2C",
		X"48",X"6E",X"72",X"6E",X"6E",X"64",X"56",X"56",X"6E",X"8B",X"77",X"51",X"35",X"19",X"3F",X"60",
		X"82",X"90",X"6E",X"4D",X"2C",X"2C",X"35",X"35",X"43",X"51",X"51",X"3A",X"1E",X"3A",X"64",X"80",
		X"A3",X"AC",X"90",X"72",X"48",X"4D",X"6E",X"90",X"B6",X"9E",X"82",X"5B",X"43",X"60",X"7C",X"A7",
		X"B1",X"90",X"77",X"48",X"4D",X"6E",X"8B",X"B6",X"A3",X"87",X"60",X"43",X"5B",X"80",X"90",X"87",
		X"8B",X"82",X"80",X"87",X"99",X"9E",X"87",X"6E",X"6E",X"95",X"B6",X"A3",X"A7",X"A3",X"95",X"80",
		X"69",X"87",X"A7",X"B6",X"95",X"72",X"4D",X"4D",X"72",X"95",X"B6",X"A7",X"82",X"60",X"43",X"27",
		X"48",X"69",X"87",X"99",X"77",X"56",X"51",X"72",X"99",X"B6",X"D7",X"CD",X"A3",X"87",X"64",X"4D",
		X"60",X"82",X"A3",X"B6",X"95",X"77",X"56",X"51",X"72",X"8B",X"B1",X"A7",X"87",X"69",X"4D",X"60",
		X"80",X"99",X"C4",X"DB",X"D2",X"BA",X"8B",X"87",X"A7",X"C8",X"D7",X"BF",X"A3",X"80",X"5B",X"72",
		X"8B",X"B6",X"CD",X"B1",X"8B",X"7C",X"95",X"BA",X"C4",X"95",X"9E",X"9E",X"99",X"A7",X"9E",X"A3",
		X"9E",X"95",X"99",X"9E",X"B1",X"BA",X"A7",X"90",X"64",X"64",X"80",X"A3",X"B6",X"A3",X"87",X"64",
		X"43",X"5B",X"77",X"9E",X"B1",X"99",X"77",X"69",X"82",X"A3",X"B6",X"B1",X"A3",X"82",X"64",X"3F",
		X"4D",X"72",X"99",X"AC",X"95",X"72",X"4D",X"3F",X"5B",X"87",X"87",X"69",X"48",X"1E",X"31",X"4D",
		X"77",X"95",X"80",X"64",X"3A",X"27",X"43",X"64",X"87",X"AC",X"B6",X"90",X"6E",X"48",X"51",X"72",
		X"69",X"6E",X"6E",X"60",X"4D",X"60",X"6E",X"64",X"6E",X"7C",X"82",X"72",X"51",X"56",X"60",X"43",
		X"2C",X"31",X"60",X"7C",X"6E",X"72",X"6E",X"5B",X"51",X"60",X"82",X"87",X"69",X"4D",X"22",X"2C",
		X"4D",X"72",X"95",X"80",X"69",X"3A",X"27",X"3A",X"31",X"3F",X"4D",X"56",X"4D",X"27",X"27",X"4D",
		X"6E",X"95",X"B1",X"A7",X"82",X"60",X"43",X"5B",X"80",X"A3",X"B6",X"99",X"72",X"4D",X"48",X"6E",
		X"90",X"B1",X"AC",X"87",X"64",X"48",X"56",X"80",X"A3",X"B6",X"9E",X"7C",X"51",X"4D",X"69",X"95",
		X"8B",X"8B",X"8B",X"80",X"82",X"8B",X"9E",X"99",X"80",X"69",X"80",X"A7",X"B1",X"A3",X"AC",X"9E",
		X"90",X"72",X"72",X"90",X"B6",X"AC",X"82",X"69",X"43",X"60",X"82",X"A3",X"BA",X"95",X"77",X"5B",
		X"35",X"31",X"56",X"72",X"95",X"90",X"6E",X"4D",X"60",X"87",X"A3",X"C4",X"D7",X"BF",X"99",X"77",
		X"51",X"4D",X"72",X"95",X"B6",X"AC",X"87",X"64",X"48",X"5B",X"82",X"A7",X"BA",X"9E",X"7C",X"56",
		X"4D",X"6E",X"90",X"B1",X"D2",X"DB",X"C8",X"A7",X"82",X"95",X"BF",X"D7",X"D2",X"B1",X"90",X"6E",
		X"60",X"82",X"9E",X"C4",X"C4",X"99",X"80",X"82",X"A7",X"C8",X"B1",X"95",X"A3",X"99",X"A3",X"A7",
		X"A3",X"A3",X"99",X"99",X"9E",X"A3",X"B6",X"B6",X"99",X"80",X"60",X"72",X"95",X"B1",X"B6",X"95",
		X"77",X"51",X"43",X"6E",X"87",X"AC",X"AC",X"82",X"64",X"6E",X"90",X"B1",X"B1",X"B1",X"95",X"72",
		X"51",X"3A",X"64",X"80",X"A3",X"A7",X"82",X"64",X"3F",X"48",X"72",X"8B",X"80",X"5B",X"35",X"22",
		X"3A",X"60",X"87",X"90",X"77",X"51",X"2C",X"2C",X"51",X"77",X"95",X"B6",X"A7",X"80",X"64",X"43",
		X"69",X"77",X"69",X"72",X"69",X"56",X"51",X"64",X"69",X"69",X"72",X"82",X"80",X"69",X"51",X"5B",
		X"56",X"3A",X"27",X"43",X"72",X"77",X"6E",X"72",X"69",X"56",X"56",X"6E",X"8B",X"82",X"60",X"3A",
		X"1E",X"35",X"60",X"82",X"95",X"77",X"56",X"2C",X"31",X"3A",X"35",X"43",X"56",X"51",X"3F",X"22",
		X"3A",X"60",X"7C",X"A3",X"B1",X"95",X"77",X"51",X"4D",X"72",X"8B",X"B1",X"A7",X"87",X"69",X"48",
		X"5B",X"80",X"9E",X"B6",X"99",X"7C",X"56",X"4D",X"6E",X"87",X"AC",X"AC",X"8B",X"6E",X"4D",X"5B",
		X"80",X"95",X"8B",X"90",X"87",X"80",X"87",X"99",X"9E",X"90",X"6E",X"6E",X"90",X"AC",X"A7",X"A7",
		X"A7",X"99",X"82",X"69",X"80",X"A7",X"BA",X"99",X"80",X"51",X"4D",X"6E",X"8B",X"B6",X"AC",X"8B",
		X"69",X"43",X"2C",X"3F",X"64",X"8B",X"99",X"82",X"5B",X"51",X"72",X"90",X"B6",X"D7",X"D7",X"AC",
		X"87",X"69",X"48",X"60",X"82",X"9E",X"BA",X"99",X"7C",X"5B",X"48",X"48",X"43",X"43",X"4D",X"56",
		X"56",X"4D",X"51",X"60",X"56",X"4D",X"5B",X"60",X"5B",X"4D",X"43",X"56",X"6E",X"90",X"BA",X"B1",
		X"90",X"72",X"4D",X"60",X"7C",X"A3",X"BF",X"A3",X"82",X"6E",X"8B",X"95",X"87",X"A3",X"9E",X"90",
		X"72",X"77",X"95",X"B6",X"AC",X"80",X"6E",X"77",X"77",X"77",X"72",X"6E",X"77",X"77",X"72",X"72",
		X"7C",X"80",X"90",X"90",X"7C",X"60",X"3A",X"51",X"77",X"95",X"AC",X"8B",X"72",X"4D",X"48",X"69",
		X"87",X"A7",X"A3",X"82",X"64",X"43",X"56",X"77",X"95",X"B1",X"95",X"77",X"56",X"48",X"69",X"87",
		X"A7",X"AC",X"87",X"6E",X"48",X"22",X"3A",X"56",X"82",X"99",X"82",X"60",X"4D",X"6E",X"87",X"AC",
		X"B6",X"90",X"77",X"51",X"5B",X"7C",X"99",X"BA",X"A7",X"87",X"64",X"4D",X"69",X"8B",X"9E",X"77",
		X"72",X"95",X"95",X"6E",X"7C",X"95",X"BA",X"DB",X"C8",X"A3",X"87",X"9E",X"BF",X"E0",X"F3",X"CD",
		X"B1",X"87",X"82",X"A3",X"C8",X"C4",X"99",X"7C",X"5B",X"3F",X"51",X"72",X"8B",X"72",X"60",X"72",
		X"5B",X"5B",X"69",X"87",X"8B",X"64",X"6E",X"72",X"56",X"3A",X"4D",X"72",X"87",X"77",X"51",X"3F",
		X"60",X"82",X"9E",X"C4",X"C4",X"A3",X"82",X"64",X"69",X"8B",X"AC",X"99",X"72",X"56",X"35",X"22",
		X"3F",X"60",X"82",X"8B",X"72",X"4D",X"48",X"72",X"90",X"B6",X"A7",X"80",X"64",X"77",X"69",X"5B",
		X"6E",X"7C",X"64",X"60",X"72",X"87",X"B6",X"AC",X"90",X"6E",X"77",X"95",X"87",X"90",X"A3",X"90",
		X"82",X"56",X"48",X"64",X"87",X"90",X"87",X"90",X"80",X"72",X"51",X"35",X"43",X"69",X"82",X"6E",
		X"48",X"3A",X"51",X"7C",X"99",X"BA",X"C4",X"99",X"80",X"5B",X"64",X"87",X"A3",X"95",X"7C",X"8B",
		X"AC",X"C8",X"A3",X"90",X"B6",X"BF",X"95",X"90",X"B6",X"B6",X"8B",X"72",X"77",X"99",X"BF",X"E0",
		X"FC",X"DB",X"B6",X"95",X"80",X"A3",X"BF",X"E5",X"E9",X"BF",X"9E",X"9E",X"C4",X"B6",X"BA",X"CD",
		X"C4",X"A3",X"90",X"A3",X"CD",X"D7",X"BA",X"95",X"90",X"95",X"8B",X"90",X"87",X"8B",X"90",X"8B",
		X"82",X"8B",X"8B",X"9E",X"A7",X"99",X"82",X"56",X"51",X"72",X"90",X"BA",X"B1",X"90",X"72",X"48",
		X"60",X"7C",X"A3",X"BF",X"9E",X"82",X"56",X"4D",X"6E",X"87",X"B6",X"B1",X"90",X"72",X"48",X"56",
		X"77",X"99",X"BA",X"9E",X"82",X"5B",X"35",X"27",X"43",X"6E",X"90",X"95",X"77",X"4D",X"56",X"77",
		X"95",X"BA",X"A3",X"87",X"60",X"48",X"64",X"80",X"AC",X"B6",X"95",X"77",X"4D",X"4D",X"6E",X"90",
		X"87",X"69",X"77",X"90",X"80",X"64",X"7C",X"9E",X"C4",X"C8",X"AC",X"80",X"7C",X"99",X"B6",X"C8",
		X"B1",X"95",X"6E",X"51",X"60",X"87",X"9E",X"82",X"69",X"3F",X"1E",X"14",X"35",X"60",X"60",X"3A",
		X"43",X"43",X"31",X"3A",X"51",X"72",X"56",X"43",X"51",X"48",X"27",X"1E",X"43",X"69",X"6E",X"4D",
		X"22",X"2C",X"51",X"72",X"99",X"B1",X"A3",X"7C",X"56",X"43",X"5B",X"87",X"90",X"77",X"56",X"2C",
		X"0B",X"10",X"35",X"60",X"80",X"72",X"4D",X"31",X"4D",X"69",X"95",X"A3",X"82",X"64",X"5B",X"69",
		X"4D",X"51",X"69",X"64",X"51",X"56",X"6E",X"8B",X"AC",X"90",X"6E",X"5B",X"77",X"82",X"7C",X"90",
		X"90",X"80",X"64",X"3F",X"48",X"72",X"8B",X"80",X"82",X"82",X"72",X"64",X"35",X"2C",X"48",X"6E",
		X"77",X"5B",X"35",X"35",X"60",X"80",X"9E",X"BA",X"AC",X"8B",X"69",X"51",X"6E",X"8B",X"A3",X"7C",
		X"77",X"90",X"B1",X"B6",X"90",X"95",X"B6",X"AC",X"87",X"99",X"B6",X"A3",X"80",X"69",X"87",X"A7",
		X"C4",X"E9",X"EE",X"C8",X"AC",X"87",X"87",X"AC",X"C8",X"E9",X"D7",X"B1",X"90",X"B1",X"C4",X"AC",
		X"C4",X"C4",X"B6",X"95",X"90",X"B6",X"D2",X"D2",X"A7",X"82",X"90",X"8B",X"90",X"8B",X"82",X"8B",
		X"8B",X"87",X"82",X"8B",X"90",X"A3",X"A3",X"8B",X"72",X"4D",X"60",X"82",X"A3",X"BF",X"9E",X"80",
		X"5B",X"48",X"72",X"8B",X"B1",X"B6",X"8B",X"6E",X"48",X"56",X"7C",X"99",X"BA",X"9E",X"7C",X"5B",
		X"43",X"69",X"82",X"A7",X"B1",X"8B",X"6E",X"4D",X"2C",X"35",X"56",X"77",X"95",X"82",X"64",X"48",
		X"64",X"87",X"A7",X"BA",X"90",X"77",X"51",X"4D",X"77",X"90",X"B6",X"A7",X"82",X"64",X"43",X"60",
		X"82",X"95",X"7C",X"69",X"87",X"95",X"72",X"6E",X"8B",X"AC",X"C4",X"B6",X"95",X"72",X"82",X"AC",
		X"BF",X"BF",X"9E",X"80",X"5B",X"4D",X"72",X"95",X"99",X"77",X"51",X"31",X"10",X"1E",X"48",X"64",
		X"51",X"3A",X"48",X"3A",X"31",X"3F",X"60",X"6E",X"48",X"48",X"4D",X"3A",X"22",X"27",X"4D",X"6E",
		X"60",X"35",X"22",X"35",X"64",X"80",X"A3",X"B1",X"8B",X"6E",X"48",X"4D",X"72",X"90",X"8B",X"64",
		X"43",X"22",X"06",X"22",X"48",X"6E",X"80",X"60",X"3A",X"35",X"56",X"7C",X"9E",X"99",X"77",X"56",
		X"64",X"60",X"4D",X"5B",X"69",X"60",X"51",X"60",X"77",X"9E",X"A3",X"82",X"64",X"69",X"8B",X"80",
		X"82",X"95",X"87",X"7C",X"4D",X"3F",X"56",X"80",X"87",X"80",X"87",X"7C",X"6E",X"4D",X"2C",X"35",
		X"60",X"7C",X"72",X"43",X"2C",X"48",X"69",X"8B",X"B6",X"BF",X"9E",X"7C",X"56",X"56",X"7C",X"9E",
		X"95",X"72",X"82",X"A7",X"BF",X"A7",X"90",X"AC",X"BA",X"9E",X"8B",X"B1",X"B6",X"95",X"6E",X"72",
		X"90",X"B1",X"DB",X"F3",X"E5",X"BA",X"90",X"80",X"95",X"BA",X"E0",X"E9",X"C8",X"9E",X"99",X"BF",
		X"B6",X"B6",X"C8",X"C4",X"A7",X"8B",X"9E",X"BF",X"D7",X"BA",X"95",X"87",X"90",X"8B",X"90",X"87",
		X"87",X"8B",X"8B",X"87",X"87",X"8B",X"95",X"A7",X"99",X"82",X"64",X"51",X"6E",X"8B",X"B1",X"B6",
		X"90",X"77",X"51",X"5B",X"7C",X"99",X"B6",X"A3",X"82",X"64",X"4D",X"69",X"82",X"A7",X"B6",X"90",
		X"77",X"51",X"51",X"77",X"90",X"B1",X"A3",X"82",X"69",X"3F",X"27",X"43",X"60",X"8B",X"95",X"7C",
		X"56",X"51",X"77",X"90",X"B6",X"AC",X"87",X"69",X"4D",X"60",X"80",X"9E",X"B6",X"99",X"7C",X"56",
		X"4D",X"6E",X"90",X"90",X"69",X"72",X"95",X"87",X"64",X"7C",X"99",X"BF",X"C4",X"AC",X"80",X"77",
		X"95",X"B6",X"C8",X"B1",X"99",X"72",X"4D",X"60",X"80",X"99",X"87",X"64",X"4D",X"1E",X"14",X"31",
		X"56",X"64",X"3F",X"43",X"48",X"31",X"3A",X"4D",X"6E",X"5B",X"3F",X"51",X"48",X"2C",X"1E",X"35",
		X"64",X"6E",X"51",X"2C",X"2C",X"51",X"6E",X"90",X"B6",X"A3",X"87",X"60",X"43",X"5B",X"80",X"90",
		X"77",X"56",X"3A",X"10",X"10",X"35",X"56",X"80",X"72",X"56",X"35",X"48",X"69",X"8B",X"A3",X"8B",
		X"69",X"56",X"69",X"51",X"4D",X"64",X"69",X"51",X"56",X"69",X"8B",X"AC",X"9E",X"77",X"5B",X"77",
		X"8B",X"7C",X"8B",X"95",X"82",X"69",X"43",X"43",X"69",X"8B",X"82",X"82",X"82",X"77",X"64",X"3F",
		X"2C",X"43",X"6E",X"7C",X"5B",X"3A",X"35",X"56",X"80",X"99",X"BF",X"B6",X"8B",X"72",X"51",X"69",
		X"8B",X"9E",X"90",X"9E",X"B6",X"DB",X"E5",X"BA",X"9E",X"7C",X"7C",X"A3",X"BF",X"E0",X"CD",X"A3",
		X"8B",X"9E",X"C8",X"DB",X"B6",X"A7",X"B1",X"AC",X"B6",X"B6",X"B1",X"B1",X"A7",X"A7",X"B1",X"BA",
		X"C8",X"BA",X"A3",X"80",X"69",X"8B",X"A7",X"CD",X"D2",X"AC",X"90",X"6E",X"72",X"90",X"B1",X"CD",
		X"BA",X"95",X"80",X"95",X"BA",X"D2",X"CD",X"C4",X"A3",X"82",X"64",X"64",X"82",X"A3",X"C4",X"B1",
		X"90",X"72",X"56",X"6E",X"90",X"A3",X"82",X"64",X"3F",X"35",X"60",X"7C",X"A3",X"99",X"77",X"56",
		X"35",X"48",X"72",X"8B",X"AC",X"C4",X"A7",X"87",X"64",X"56",X"80",X"7C",X"77",X"7C",X"6E",X"5B",
		X"64",X"77",X"6E",X"72",X"82",X"8B",X"82",X"69",X"5B",X"64",X"56",X"3A",X"35",X"5B",X"7C",X"77",
		X"77",X"77",X"69",X"5B",X"60",X"7C",X"90",X"77",X"56",X"35",X"22",X"4D",X"69",X"90",X"90",X"69",
		X"4D",X"2C",X"35",X"35",X"3A",X"4D",X"56",X"51",X"35",X"22",X"48",X"69",X"87",X"AC",X"AC",X"8B",
		X"6E",X"4D",X"56",X"77",X"95",X"B1",X"9E",X"80",X"5B",X"48",X"64",X"82",X"A7",X"AC",X"8B",X"72",
		X"4D",X"51",X"77",X"90",X"B1",X"9E",X"82",X"60",X"48",X"60",X"82",X"90",X"87",X"8B",X"80",X"80",
		X"8B",X"99",X"99",X"82",X"64",X"72",X"95",X"AC",X"A3",X"A7",X"9E",X"90",X"77",X"69",X"82",X"AC",
		X"AC",X"8B",X"6E",X"43",X"51",X"77",X"9E",X"B1",X"A3",X"7C",X"56",X"35",X"22",X"4D",X"69",X"90",
		X"95",X"6E",X"4D",X"51",X"7C",X"99",X"BA",X"D7",X"BF",X"99",X"80",X"5B",X"48",X"69",X"82",X"A7",
		X"AC",X"8B",X"72",X"4D",X"51",X"77",X"95",X"B1",X"9E",X"80",X"60",X"48",X"60",X"82",X"9E",X"C8",
		X"DB",X"CD",X"B1",X"82",X"8B",X"A7",X"C8",X"D2",X"B6",X"99",X"72",X"56",X"77",X"90",X"BA",X"C4",
		X"A7",X"82",X"7C",X"99",X"BF",X"BA",X"90",X"9E",X"95",X"9E",X"A3",X"9E",X"9E",X"99",X"95",X"99",
		X"9E",X"B1",X"B6",X"A3",X"87",X"5B",X"69",X"82",X"A3",X"B6",X"9E",X"80",X"56",X"3F",X"60",X"77",
		X"A3",X"AC",X"90",X"6E",X"69",X"87",X"A7",X"B1",X"AC",X"99",X"7C",X"56",X"3A",X"56",X"72",X"99",
		X"AC",X"8B",X"72",X"43",X"3F",X"60",X"82",X"82",X"60",X"43",X"22",X"31",X"56",X"77",X"90",X"77",
		X"5B",X"35",X"27",X"48",X"69",X"87",X"B1",X"AC",X"8B",X"69",X"43",X"56",X"72",X"69",X"6E",X"69",
		X"5B",X"4D",X"60",X"69",X"60",X"6E",X"7C",X"82",X"6E",X"4D",X"56",X"5B",X"3F",X"22",X"35",X"60",
		X"72",X"69",X"6E",X"69",X"56",X"51",X"64",X"87",X"82",X"64",X"43",X"19",X"31",X"51",X"77",X"95",
		X"77",X"60",X"31",X"27",X"35",X"31",X"3F",X"51",X"56",X"43",X"22",X"2C",X"51",X"72",X"99",X"B1",
		X"9E",X"7C",X"56",X"43",X"60",X"82",X"A7",X"B1",X"90",X"69",X"48",X"4D",X"72",X"95",X"B1",X"A3",
		X"80",X"5B",X"43",X"60",X"82",X"A7",X"B1",X"95",X"6E",X"4D",X"4D",X"6E",X"95",X"87",X"8B",X"87",
		X"80",X"82",X"90",X"9E",X"90",X"77",X"69",X"87",X"AC",X"AC",X"A3",X"A7",X"99",X"8B",X"6E",X"77",
		X"99",X"B6",X"9E",X"7C",X"60",X"43",X"69",X"82",X"A7",X"B1",X"8B",X"6E",X"51",X"2C",X"35",X"5B",
		X"7C",X"95",X"87",X"64",X"4D",X"69",X"8B",X"A7",X"CD",X"D7",X"B6",X"95",X"77",X"48",X"56",X"72",
		X"95",X"BA",X"A3",X"87",X"60",X"48",X"64",X"80",X"AC",X"B6",X"95",X"7C",X"4D",X"51",X"72",X"90",
		X"B6",X"D7",X"DB",X"C4",X"99",X"82",X"95",X"BF",X"D7",X"CD",X"B1",X"87",X"64",X"60",X"82",X"A7",
		X"C8",X"BF",X"99",X"77",X"87",X"A7",X"C4",X"A7",X"95",X"A3",X"99",X"A7",X"A3",X"A3",X"9E",X"99",
		X"99",X"9E",X"A7",X"BA",X"AC",X"95",X"77",X"5B",X"7C",X"99",X"B1",X"B1",X"8B",X"72",X"48",X"48",
		X"72",X"8B",X"B1",X"A3",X"7C",X"64",X"72",X"99",X"B6",X"B1",X"AC",X"8B",X"6E",X"48",X"3F",X"69",
		X"82",X"AC",X"A3",X"7C",X"60",X"3F",X"51",X"7C",X"8B",X"7C",X"51",X"2C",X"22",X"43",X"69",X"8B",
		X"8B",X"6E",X"48",X"27",X"31",X"5B",X"80",X"99",X"BA",X"9E",X"7C",X"5B",X"43",X"6E",X"72",X"69",
		X"72",X"64",X"51",X"51",X"69",X"64",X"69",X"77",X"82",X"80",X"60",X"51",X"5B",X"51",X"35",X"27",
		X"4D",X"77",X"72",X"6E",X"72",X"64",X"56",X"5B",X"77",X"8B",X"7C",X"56",X"31",X"1E",X"3F",X"64",
		X"87",X"90",X"72",X"4D",X"27",X"31",X"35",X"35",X"48",X"56",X"51",X"35",X"22",X"3A",X"64",X"82",
		X"A7",X"B1",X"8B",X"72",X"4D",X"4D",X"77",X"90",X"B6",X"A3",X"80",X"60",X"43",X"64",X"82",X"A3",
		X"B6",X"90",X"77",X"51",X"4D",X"77",X"90",X"B6",X"A7",X"82",X"64",X"48",X"5B",X"87",X"95",X"87",
		X"90",X"82",X"82",X"87",X"9E",X"9E",X"8B",X"72",X"72",X"95",X"B1",X"A7",X"A7",X"A3",X"95",X"7C",
		X"69",X"82",X"AC",X"B6",X"90",X"77",X"48",X"56",X"72",X"95",X"BA",X"A3",X"87",X"64",X"3A",X"27",
		X"43",X"6E",X"90",X"99",X"7C",X"51",X"56",X"77",X"95",X"BF",X"DB",X"CD",X"A3",X"82",X"64",X"48",
		X"64",X"87",X"A7",X"BA",X"90",X"77",X"51",X"4D",X"77",X"90",X"B6",X"A7",X"82",X"64",X"48",X"60",
		X"82",X"A3",X"C4",X"DB",X"D2",X"B6",X"90",X"8B",X"AC",X"CD",X"D7",X"BF",X"9E",X"80",X"60",X"72",
		X"90",X"B6",X"C8",X"AC",X"87",X"7C",X"99",X"BF",X"C4",X"99",X"9E",X"9E",X"99",X"A7",X"9E",X"A3",
		X"9E",X"99",X"99",X"9E",X"AC",X"BA",X"A7",X"8B",X"69",X"64",X"82",X"A3",X"B6",X"A3",X"82",X"64",
		X"48",X"5B",X"7C",X"9E",X"B1",X"95",X"72",X"64",X"87",X"A7",X"B6",X"B1",X"9E",X"80",X"60",X"43",
		X"51",X"72",X"90",X"AC",X"90",X"77",X"51",X"43",X"60",X"82",X"8B",X"64",X"48",X"22",X"2C",X"56",
		X"72",X"95",X"80",X"5B",X"3A",X"22",X"43",X"69",X"82",X"A7",X"B1",X"90",X"72",X"4D",X"51",X"77",
		X"6E",X"6E",X"6E",X"60",X"4D",X"60",X"6E",X"64",X"6E",X"80",X"87",X"72",X"51",X"56",X"60",X"43",
		X"27",X"35",X"60",X"77",X"6E",X"72",X"6E",X"5B",X"56",X"64",X"80",X"87",X"69",X"48",X"27",X"2C",
		X"51",X"72",X"90",X"80",X"64",X"3F",X"2C",X"3A",X"35",X"3F",X"51",X"56",X"48",X"2C",X"2C",X"51",
		X"6E",X"90",X"B6",X"A3",X"82",X"60",X"43",X"60",X"7C",X"A7",X"B6",X"95",X"77",X"4D",X"4D",X"6E",
		X"90",X"B6",X"A7",X"87",X"64",X"43",X"60",X"7C",X"A3",X"B6",X"95",X"7C",X"4D",X"4D",X"6E",X"90",
		X"8B",X"8B",X"8B",X"80",X"82",X"90",X"9E",X"95",X"7C",X"69",X"7C",X"A7",X"B1",X"A3",X"AC",X"99",
		X"90",X"6E",X"72",X"99",X"B6",X"AC",X"82",X"60",X"48",X"60",X"82",X"A7",X"B6",X"99",X"72",X"56",
		X"31",X"31",X"5B",X"77",X"99",X"90",X"69",X"4D",X"60",X"87",X"A7",X"C8",X"DB",X"BA",X"95",X"7C",
		X"56",X"51",X"72",X"90",X"B1",X"AC",X"87",X"69",X"48",X"48",X"48",X"48",X"95",X"A7",X"9E",X"A3",
		X"9E",X"9E",X"9E",X"9E",X"9E",X"9E",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"95",X"95",X"95",
		X"95",X"95",X"95",X"95",X"95",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"8B",X"8B",
		X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"8B",X"87",X"87",X"87",X"87",X"87",X"87",X"87",
		X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"87",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",
		X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"82",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",
		X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C",X"7C");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
